module prod
(
  input clk, 
);

//(* gclk *) wire clk;

//**Wire declarations**//
//**Init register**//
//**Stuttering Signal**//
//**Self-composed modules**//
//**Initial state**//
//**State invariants**//
//**Verification conditions**//

endmodule