module SodorInternalTile_1stage_inductive_state_src ( input \Core_1stage.DatPath_1stage.reg_interrupt_edge , input [31:0] \Core_1stage.DatPath_1stage.if_inst_buffer , input \Core_1stage.CtlPath_1stage.reg_mem_en , input \Core_1stage.DatPath_1stage.reg_dmiss , output \Core_1stage.CtlPath_1stage.reg_mem_en_inductive_state_src , output \Core_1stage.DatPath_1stage.reg_dmiss_inductive_state_src , output [31:0] \Core_1stage.DatPath_1stage.if_inst_buffer_inductive_state_src , output \Core_1stage.DatPath_1stage.reg_interrupt_edge_inductive_state_src );
	assign \Core_1stage.DatPath_1stage.reg_dmiss_inductive_state_src = \Core_1stage.DatPath_1stage.reg_dmiss ;
	assign \Core_1stage.DatPath_1stage.if_inst_buffer_inductive_state_src = \Core_1stage.DatPath_1stage.if_inst_buffer ;
	assign \Core_1stage.DatPath_1stage.reg_interrupt_edge_inductive_state_src = \Core_1stage.DatPath_1stage.reg_interrupt_edge ;
	assign \Core_1stage.CtlPath_1stage.reg_mem_en_inductive_state_src = \Core_1stage.CtlPath_1stage.reg_mem_en ;
endmodule