module SodorInternalTile_2stage_obs_trg ( input \Core_2stage.c_io_dat_mem_store , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_192 , input \Core_2stage.DatPath_2stage._exe_wbdata_T_2 , input [6:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_2 , input [4:0] \Core_2stage.DatPath_2stage.alu_shamt , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_127 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_183 , input [31:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data , input \Core_2stage.io_interrupt_msip , input [9:0] \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_addr , input [4:0] \Core_2stage.DatPath_2stage.exe_rs2_addr , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_617 , input \Core_2stage.DatPath_2stage._exe_alu_op2_T_3 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_wfi , input [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_0 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_3 , input \Core_2stage.DatPath_2stage._csr_io_tval_T_2 , input [31:0] \Core_2stage.DatPath_2stage.imm_z , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_3 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_3 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_226 , input core_io_interrupt_meip , input [31:0] router_1_io_corePort_req_bits_addr , input \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugBreak , input [2:0] \Core_2stage.CtlPath_2stage.io_dmem_req_bits_typ , input \Core_2stage.DatPath_2stage._if_pc_next_T_4 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_364 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_376 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_26 , input [2:0] \Core_2stage.CtlPath_2stage.io_ctl_mem_typ , input \Core_2stage.d_io_interrupt_debug , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_3 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_172 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_3 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_34 , input [31:0] router_io_corePort_req_bits_data , input \Core_2stage.CtlPath_2stage._csignals_T_5 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_335 , input \SodorRequestRouter_2stage_0.in_range , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_117 , input [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_cmd , input \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_0 , input [9:0] \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_addr , input [32:0] \SodorRequestRouter_2stage_1._in_range_T_1 , input [31:0] io_debug_port_resp_bits_data , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_31 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._notDebugTVec_T_1 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_23 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_322 , input \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_signed , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_11 , input \Core_2stage.CtlPath_2stage._csignals_T_95 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_26 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_13 , input [31:0] io_master_port_1_resp_bits_data , input \Core_2stage.DatPath_2stage._exe_alu_out_T_21 , input [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_1 , input [31:0] \Core_2stage.DatPath_2stage.regfile_14 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_121 , input [2:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_req_bits_typ , input \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_2 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_316 , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._bytes_T_1 , input \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_mask , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_mtip , input [7:0] \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_data , input \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_signed_state_invariant , input [31:0] \Core_2stage.DatPath_2stage.regfile_1 , input \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_en , input [2:0] \SodorRequestRouter_2stage_1.io_corePort_req_bits_typ , input [7:0] \Core_2stage.DatPath_2stage._T_17 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.new_dcsr_ebreakm , input [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._large_r_T_1 , input \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_en , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_size , input [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_24 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_324 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_1 , input [31:0] \Core_2stage.DatPath_2stage.regfile_23 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_312 , input [31:0] \Core_2stage.DatPath_2stage.exe_wbdata , input \Core_2stage.DatPath_2stage._exe_alu_out_T_25 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_2 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_238 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_9 , input \Core_2stage.DatPath_2stage.csr_io_status_upie , input \Core_2stage.DatPath_2stage.CSRFile_2stage._T_15 , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_3 , input [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_170 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_193 , input \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_1 , input [1:0] \Core_2stage.c_io_ctl_op1_sel , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_618 , input [9:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_addr , input [2:0] router_io_masterPort_req_bits_typ , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mscratch , input \Core_2stage.DatPath_2stage.csr_io_status_tvm , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_12 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_upie , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_119 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_306 , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_3 , input \Core_2stage.d_io_ctl_stall , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_hie , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_627 , input [2:0] \AsyncScratchPadMemory_2stage._io_core_ports_1_resp_bits_data_T_1 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_637 , input \Core_2stage.CtlPath_2stage._csignals_T_87 , input [31:0] io_master_port_0_req_bits_addr , input [10:0] \Core_2stage.DatPath_2stage._imm_j_sext_T_2 , input \Core_2stage.d_io_imem_req_valid , input [7:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.cause_lsbs , input [31:0] \Core_2stage.DatPath_2stage.io_dmem_resp_bits_data , input [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_2 , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_316 , input io_interrupt_msip , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_195 , input [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_mask , input [31:0] core_io_imem_req_bits_addr , input [31:0] \Core_2stage.io_imem_resp_bits_data_state_invariant , input [31:0] \Core_2stage.DatPath_2stage.regfile_15 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._epc_T_1 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dpc , input \Core_2stage.CtlPath_2stage.io_dat_data_misaligned , input \Core_2stage.d_io_dat_br_eq , input \Core_2stage.d_io_interrupt_msip , input [8:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_lo_lo , input [31:0] router_io_respAddress , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_4 , input \Core_2stage.DatPath_2stage._exe_wbdata_T_3 , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._bytes_T_3 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_586 , input [5:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.small_ , input \Core_2stage.DatPath_2stage.CSRFile_2stage._io_eret_T , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_14 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mbe , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_206 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_383 , input router_1_io_masterPort_req_valid , input [5:0] \Core_2stage.DatPath_2stage._misaligned_mask_T_3 , input \Core_2stage.c_io_ctl_rf_wen , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_123 , input [2:0] io_debug_port_req_bits_typ , input [31:0] io_debug_port_req_bits_addr , input \Core_2stage.DatPath_2stage.csr_io_eret , input [31:0] \Core_2stage.DatPath_2stage.regfile_25 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_285 , input [62:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_19 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_359 , input [31:0] \SodorRequestRouter_2stage_1.io_corePort_req_bits_data , input \Core_2stage.DatPath_2stage.io_ctl_if_kill_r , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_27 , input \Core_2stage.CtlPath_2stage._csignals_T_63 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_175 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.new_mstatus_mpie , input [31:0] core_io_dmem_req_bits_data , input [7:0] \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_data , input [31:0] router_io_masterPort_resp_bits_data , input [7:0] \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_data , input [1:0] \Core_2stage.d_io_ctl_op1_sel , input core_io_imem_req_valid , input [7:0] \AsyncScratchPadMemory_2stage.module_1_io_mem_data_1 , input \AsyncScratchPadMemory_2stage.module__io_en , input [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data , input [31:0] \Core_2stage.DatPath_2stage.io_ctl_exception_cause , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_3 , input [31:0] \Core_2stage.d_io_imem_req_bits_addr , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_293 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_18 , input [31:0] \Core_2stage.DatPath_2stage.if_reg_pc , input [31:0] \Core_2stage.DatPath_2stage.regfile_18 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_393 , input \Core_2stage.DatPath_2stage.io_dat_data_misaligned , input [2:0] \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_1 , input \Core_2stage.DatPath_2stage.reg_interrupt_handled , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_2 , input [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.large_1 , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.value_1 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_3 , input [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.offset , input core_io_dmem_req_bits_fcn , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_217 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._epc_T , input [31:0] \Core_2stage.DatPath_2stage.exception_target , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_373 , input [31:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_data , input [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.large_ , input \Core_2stage.DatPath_2stage.io_dat_mem_store , input clock , input [4:0] \Core_2stage.c_io_ctl_alu_fun , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_2 , input [31:0] \AsyncScratchPadMemory_2stage.module__io_data , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_msip , input [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_3 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_19 , input \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_2 , input [10:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._masks_mask_T , input \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_0 , input [7:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_2 , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_en , input \Core_2stage.CtlPath_2stage._csignals_T_97 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_35 , input [31:0] \Core_2stage.DatPath_2stage.io_reset_vector , input \Core_2stage.DatPath_2stage.csr_io_retire , input \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_13 , input \Core_2stage.d_io_ctl_rf_wen , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_184 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_11 , input [7:0] \Core_2stage.DatPath_2stage._T_6 , input [2:0] \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_typ , input [9:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_addr , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.s_offset , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_3 , input [31:0] \Core_2stage.DatPath_2stage.csr_io_interrupt_cause , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_1 , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_20 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_retire , input [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_size , input [7:0] \AsyncScratchPadMemory_2stage.mem_2_MPORT_data , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_5 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_7 , input [9:0] \AsyncScratchPadMemory_2stage.module__io_mem_addr , input [31:0] \Core_2stage.DatPath_2stage.regfile_4 , input [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_5 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sum , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_185 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_179 , input [20:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_addr , input \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_1 , input \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_valid , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_246 , input [2:0] \Core_2stage.d_io_ctl_mem_typ , input [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_21 , input reset , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_interruptVec , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_622 , input [31:0] \Core_2stage.d_io_ctl_exception_cause , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_10 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_debug , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_31 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_3 , input [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._large_r_T_3 , input io_master_port_1_req_bits_fcn , input \Core_2stage.DatPath_2stage._if_pc_next_T_3 , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_mask , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_274 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_2 , input [31:0] \Core_2stage.DatPath_2stage._if_pc_next_T_6 , input [7:0] \AsyncScratchPadMemory_2stage.module_1_io_mem_data_2 , input [7:0] \Core_2stage.DatPath_2stage._T_8 , input \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_274 , input [31:0] \Core_2stage.DatPath_2stage.if_inst_buffer , input \Core_2stage.CtlPath_2stage._csignals_T_71 , input \Core_2stage.DatPath_2stage.io_dat_br_ltu , input core_io_interrupt_mtip , input router_1_io_corePort_req_valid , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_284 , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_115 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_295 , input \Core_2stage.d_io_dat_csr_eret , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_10 , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_123 , input [31:0] \Core_2stage.DatPath_2stage.regfile_3 , input \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_273 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_meip , input \AsyncScratchPadMemory_2stage.MemReader_2stage_2.sign , input \Core_2stage.DatPath_2stage.csr_io_interrupts_debug , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_363 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_281 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_245 , input [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_8 , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_109 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_18 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugInt , input [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_30 , input [2:0] \Core_2stage.DatPath_2stage.io_ctl_csr_cmd , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_178 , input \Core_2stage.CtlPath_2stage._csignals_T_436 , input [31:0] \Core_2stage.DatPath_2stage.regfile_MPORT_data , input [1:0] \Core_2stage.DatPath_2stage.csr_io_status_sxl , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_344 , input \Core_2stage.DatPath_2stage.io_imem_req_valid , input [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_hi , input [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_cause , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_619 , input \AsyncScratchPadMemory_2stage.io_debug_port_req_valid , input [62:0] \Core_2stage.DatPath_2stage._GEN_11 , input \Core_2stage.DatPath_2stage.csr_io_status_sbe , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_286 , input [15:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mip , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_126 , input router_1_io_masterPort_req_bits_fcn , input [4:0] \Core_2stage.CtlPath_2stage.io_ctl_alu_fun , input \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_3 , input \Core_2stage.d_io_dat_data_misaligned , input [1:0] \Core_2stage.DatPath_2stage.csr_io_status_mpp , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_280 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_debug , input \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_en , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_mask , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_2 , input [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_2 , input [31:0] \Core_2stage.d_io_dmem_req_bits_data , input \Core_2stage.io_interrupt_meip , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_370 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_602 , input [31:0] \Core_2stage.DatPath_2stage.csr_io_rw_rdata , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_610 , input [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_1 , input \SodorRequestRouter_2stage_0.io_masterPort_req_bits_fcn , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mcountinhibit_T_1 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_op2_T_6 , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugBreak_T_4 , input [18:0] \Core_2stage.DatPath_2stage._imm_b_sext_T_2 , input router_1_io_corePort_req_bits_fcn , input \Core_2stage.DatPath_2stage._exe_alu_op2_T_1 , input [32:0] \SodorRequestRouter_2stage_1._resp_in_range_T_1 , input [4:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._shiftedVec_T , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_187 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_5 , input \Core_2stage.c_io_dmem_resp_valid , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_spp , input [2:0] \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_typ , input \Core_2stage.CtlPath_2stage._csignals_T_85 , input \Core_2stage.CtlPath_2stage._csignals_T_79 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_isa , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_10 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_3 , input [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_5 , input [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_size , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_20 , input \Core_2stage.CtlPath_2stage._csignals_T_1 , input \Core_2stage.DatPath_2stage._exe_alu_out_T_8 , input \SodorRequestRouter_2stage_1.io_masterPort_req_bits_fcn , input \Core_2stage.CtlPath_2stage._csignals_T_49 , input \Core_2stage.CtlPath_2stage.io_ctl_exception , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_3 , input [7:0] \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_data , input [6:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_maskWithOffset_T , input [7:0] \AsyncScratchPadMemory_2stage.mem_1_MPORT_data , input \Core_2stage.d_io_interrupt_meip , input [31:0] \Core_2stage.DatPath_2stage.csr_io_cause , input [20:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_addr_state_invariant , input [7:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_3 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_2 , input [2:0] core_io_dmem_req_bits_typ , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_219 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_243 , input \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_en , input [104:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._new_mstatus_WIRE , input router_io_masterPort_req_bits_fcn , input \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_wfi , input [7:0] \AsyncScratchPadMemory_2stage.module_1_io_mem_data_0 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_368 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_625 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_353 , input [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_dprv , input [2:0] io_master_port_1_req_bits_typ , input [2:0] memory_io_core_ports_1_req_bits_typ , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_292 , input [31:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_data , input [19:0] \Core_2stage.DatPath_2stage._imm_i_sext_T_2 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_611 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_181 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_229 , input [2:0] \Core_2stage.CtlPath_2stage.cs0_4 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_176 , input [7:0] \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_data , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupt , input core_io_imem_resp_valid , input \Core_2stage.DatPath_2stage.io_ctl_mem_val , input [10:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._masks_mask_T , input \Core_2stage.CtlPath_2stage._csignals_T_33 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_309 , input \Core_2stage.DatPath_2stage._exe_alu_op1_T_2 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_dv , input [2:0] \Core_2stage.CtlPath_2stage.csr_cmd , input \Core_2stage.CtlPath_2stage._csignals_T_27 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_342 , input [11:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_addr , input \SodorRequestRouter_2stage_0.io_masterPort_req_valid , input [31:0] \SodorRequestRouter_2stage_1.io_corePort_resp_bits_data , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_3 , input \SodorRequestRouter_2stage_0.resp_in_range , input \Core_2stage.c_io_dat_csr_interrupt , input \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_2 , input [9:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_addr_state_invariant , input \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_signed , input [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_uxl , input [31:0] router_1_io_scratchPort_req_bits_addr , input [22:0] \Core_2stage.DatPath_2stage.csr_io_status_zero2 , input \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_7 , input [11:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._debugTVec_T , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpie , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_392 , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_121 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_380 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_0 , input [9:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_addr , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_365 , input \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_signed , input [31:0] \Core_2stage.d_io_reset_vector , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_3 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_221 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_116 , input \Core_2stage.DatPath_2stage.CSRFile_2stage._T_183 , input [31:0] \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_data , input [20:0] \AsyncScratchPadMemory_2stage.module_1_io_addr , input router_1_io_scratchPort_req_bits_fcn , input [31:0] core_io_reset_vector , input \Core_2stage.DatPath_2stage.csr_io_status_mpv , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_146 , input \Core_2stage.CtlPath_2stage.io_imem_resp_valid , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_601 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_14 , input [10:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._masks_mask_T , input \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_mask , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_111 , input [31:0] \Core_2stage.c_io_ctl_exception_cause , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_358 , input [31:0] \SodorRequestRouter_2stage_1.io_respAddress , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_1 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_17 , input [31:0] memory_io_core_ports_0_resp_bits_data , input [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_maskWithOffset , input \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugTrigger , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_2 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.tvec , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo , input \Core_2stage.DatPath_2stage.csr_io_status_sum , input \Core_2stage.c_io_ctl_stall , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_16 , input [9:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_addr , input [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_3 , input [20:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_addr , input \Core_2stage.d_io_interrupt_mtip , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_1 , input \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_en , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_8 , input \Core_2stage.DatPath_2stage.csr_io_status_v , input \Core_2stage.io_interrupt_mtip , input [31:0] io_master_port_0_resp_bits_data , input [31:0] \SodorRequestRouter_2stage_0.io_masterPort_req_bits_data , input [10:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._masks_mask_T , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.pending_interrupts , input \Core_2stage.DatPath_2stage._exe_alu_out_T_27 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_15 , input \AsyncScratchPadMemory_2stage.mem_2_MPORT_en , input router_1_io_masterPort_resp_valid , input [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_0 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_307 , input \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_178 , input [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_1 , input \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_en , input [7:0] \Core_2stage.DatPath_2stage._T_5 , input \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_11 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_28 , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_346 , input [32:0] \SodorRequestRouter_2stage_1._resp_in_range_T_3 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_13 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_196 , input \Core_2stage.CtlPath_2stage._csignals_T_11 , input [31:0] router_1_io_corePort_resp_bits_data , input \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_mask , input \Core_2stage.CtlPath_2stage._csignals_T_31 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_27 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_231 , input [7:0] \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_data , input \Core_2stage.CtlPath_2stage._csignals_T_81 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_276 , input [2:0] \Core_2stage.d_io_ctl_pc_sel , input \Core_2stage.CtlPath_2stage._csignals_T_538 , input \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_182 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_1 , input \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_12 , input [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_3 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_313 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_385 , input [31:0] router_1_io_masterPort_req_bits_data , input \Core_2stage.DatPath_2stage.CSRFile_2stage.x86 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_275 , input [31:0] \SodorRequestRouter_2stage_0.io_scratchPort_resp_bits_data , input [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_hi , input [31:0] \Core_2stage.DatPath_2stage.io_dat_inst , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_ebreakm , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_spie , input [104:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mstatus_T , input \Core_2stage.c_io_ctl_exception , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_3 , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_294 , input \Core_2stage.DatPath_2stage.csr_io_exception , input [9:0] \AsyncScratchPadMemory_2stage.mem_1_MPORT_addr , input \SodorRequestRouter_2stage_0.io_scratchPort_req_valid , input \Core_2stage.CtlPath_2stage._csignals_T_51 , input \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_2 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_615 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_587 , input [2:0] \Core_2stage.d_io_ctl_op2_sel , input [31:0] core_io_dmem_resp_bits_data , input [31:0] \Core_2stage.DatPath_2stage.io_dmem_req_bits_data , input [1:0] \Core_2stage.DatPath_2stage.csr_io_status_fs , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_3 , input memory_io_core_ports_1_resp_valid , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_106 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_215 , input \Core_2stage.DatPath_2stage._exe_alu_out_T_12 , input \AsyncScratchPadMemory_2stage.module__io_mem_masks_2 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_378 , input \SodorRequestRouter_2stage_0.io_corePort_resp_valid , input \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_1 , input [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_hi , input [7:0] \Core_2stage.DatPath_2stage._T_16 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_291 , input \Core_2stage.CtlPath_2stage._csignals_T_410 , input \Core_2stage.CtlPath_2stage._csignals_T_77 , input \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_signed , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_616 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_26 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_212 , input [7:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_0 , input \AsyncScratchPadMemory_2stage.MemReader_2stage_1.sign , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_2 , input \Core_2stage.CtlPath_2stage.io_dmem_resp_valid , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_11 , input [4:0] \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_addr , input \SodorRequestRouter_2stage_1.io_corePort_req_bits_fcn , input [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_214 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_2 , input \Core_2stage.c_io_dmem_req_bits_fcn , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_0 , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_3 , input \Core_2stage.c_io_dat_br_eq , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tw , input [31:0] \SodorRequestRouter_2stage_1.io_scratchPort_resp_bits_data , input \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_2 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_31 , input [15:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mip_T , input [21:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_lo , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_3 , input [20:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_addr , input [2:0] \Core_2stage.CtlPath_2stage.ctrl_pc_sel_no_xept , input \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_en , input \Core_2stage.CtlPath_2stage._csignals_T_55 , input [31:0] \SodorRequestRouter_2stage_1.io_masterPort_req_bits_data , input [9:0] \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_addr , input \Core_2stage.DatPath_2stage._exe_alu_out_T , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_32 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupt_cause , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_27 , input \Core_2stage.DatPath_2stage._csr_io_tval_T_3 , input [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_prv , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_15 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.trapToDebug , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_208 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_3 , input [9:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_addr , input \Core_2stage.CtlPath_2stage.cs0_2 , input [31:0] \Core_2stage.CtlPath_2stage._csignals_T_38 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_107 , input [6:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._GEN_1 , input [31:0] \Core_2stage.DatPath_2stage._exe_wbdata_T_4 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_624 , input \Core_2stage.DatPath_2stage.CSRFile_2stage._T_368 , input [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_1_state_invariant , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_236 , input [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_maskWithOffset , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_0 , input \Core_2stage.DatPath_2stage._exe_alu_op1_T , input [9:0] \AsyncScratchPadMemory_2stage.mem_2_MPORT_addr , input [82:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_hi , input \AsyncScratchPadMemory_2stage.io_debug_port_resp_valid , input [31:0] memory_io_core_ports_1_req_bits_addr , input \Core_2stage.d_io_dat_br_ltu , input \Core_2stage.DatPath_2stage.io_dat_csr_eret , input \Core_2stage.CtlPath_2stage._csignals_T_91 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_exception , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_240 , input [31:0] \Core_2stage.DatPath_2stage.regfile_19 , input [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_lo , input [9:0] \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_addr , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.s_offset , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_tval , input [7:0] \Core_2stage.DatPath_2stage._T_12 , input \AsyncScratchPadMemory_2stage.module__io_mem_masks_1 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_327 , input [4:0] \Core_2stage.DatPath_2stage.regfile_MPORT_addr , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_328 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_390 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_367 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.clock , input [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_mask , input [31:0] \Core_2stage.DatPath_2stage.csr_io_pc , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_30 , input [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data , input io_interrupt_mtip , input [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_15 , input [9:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_addr , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_119 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_315 , input [31:0] \Core_2stage.d_io_dmem_resp_bits_data , input \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_0 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_0 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_266 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_15 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_hartid , input [9:0] \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_addr , input \Core_2stage.DatPath_2stage.regfile_MPORT_1_mask , input \SodorRequestRouter_2stage_1.io_scratchPort_req_valid , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_2 , input [31:0] router_1_io_scratchPort_resp_bits_data , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._sign_T_1 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_596 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_607 , input \AsyncScratchPadMemory_2stage.MemReader_2stage_0.sign , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_37 , input [31:0] \Core_2stage.io_imem_req_bits_addr , input \SodorRequestRouter_2stage_0.io_corePort_req_valid , input \Core_2stage.DatPath_2stage.CSRFile_2stage._any_T_78 , input \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_en , input \Core_2stage.c_io_dat_if_valid_resp , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_220 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_6 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mxr , input [31:0] \Core_2stage.DatPath_2stage.regfile_11 , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_101 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_15 , input [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_mask , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mcause_T , input [6:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_interruptOffset , input [31:0] router_io_corePort_resp_bits_data , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_343 , input \Core_2stage.CtlPath_2stage.io_ctl_stall , input [31:0] \SodorRequestRouter_2stage_0.io_masterPort_req_bits_addr , input \Core_2stage.d_io_hartid , input \Core_2stage.DatPath_2stage.csr_io_status_uie , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_4 , input [7:0] \Core_2stage.DatPath_2stage.csr_io_status_zero1 , input io_master_port_0_req_valid , input [62:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._GEN_0 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_294 , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_99 , input [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_3 , input [4:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._shiftedVec_T , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_583 , input core_clock , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_621 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_24 , input \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_8 , input \AsyncScratchPadMemory_2stage.clock , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mie , input [2:0] \Core_2stage.c_io_ctl_mem_typ , input [31:0] router_io_scratchPort_req_bits_addr , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_361 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mtvec , input \Core_2stage.CtlPath_2stage._csignals_T_61 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_debug , input [31:0] io_imem_req_bits_addr_state_invariant , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_223 , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_0 , input [31:0] \Core_2stage.DatPath_2stage.exe_reg_pc_plus4 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tsr , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_22 , input [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_2 , input \Core_2stage.d_io_ctl_if_kill , input [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_maskWithOffset , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtvec , input [7:0] \Core_2stage.DatPath_2stage._T_10 , input [2:0] \Core_2stage.DatPath_2stage.io_ctl_pc_sel_no_xept , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_7 , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1722 , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_26 , input [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.offset , input [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_73 , input [31:0] \Core_2stage.DatPath_2stage.regfile_7 , input \Core_2stage.CtlPath_2stage._csignals_T_437 , input [20:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_addr , input [31:0] router_io_masterPort_req_bits_data , input \Core_2stage.DatPath_2stage.CSRFile_2stage.new_mstatus_mie , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_11 , input \AsyncScratchPadMemory_2stage.module__io_mem_masks_3 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_222 , input [7:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_1 , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_en , input [31:0] router_1_io_masterPort_resp_bits_data , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_8 , input [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_19 , input \Core_2stage.DatPath_2stage._exe_wbdata_T_1 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_321 , input [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_25 , input \Core_2stage.CtlPath_2stage._csignals_T_93 , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_345 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_23 , input [5:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_34 , input [2:0] \Core_2stage.io_dmem_req_bits_typ , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_maskWithOffset , input \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_145 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_ret , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_29 , input [31:0] \Core_2stage.DatPath_2stage.regfile_2 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_26 , input \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_217 , input \AsyncScratchPadMemory_2stage.mem_1_MPORT_mask , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._bytes_T_1 , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_1 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_break , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_227 , input \Core_2stage.c_io_dat_br_ltu , input \Core_2stage.DatPath_2stage.CSRFile_2stage._io_decode_0_read_illegal_T_16 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_23 , input \Core_2stage.c_io_dat_csr_eret , input [9:0] \AsyncScratchPadMemory_2stage.mem_3_MPORT_addr , input \Core_2stage.c_io_imem_resp_valid , input [31:0] \Core_2stage.DatPath_2stage.exe_jmp_target , input [31:0] \Core_2stage.io_dmem_resp_bits_data , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_122 , input \Core_2stage.CtlPath_2stage._csignals_T_408 , input [9:0] \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_addr , input [31:0] memory_io_core_ports_1_resp_bits_data , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_singleStep , input [22:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_zero2 , input \Core_2stage.CtlPath_2stage.io_dat_csr_interrupt , input \Core_2stage.d_io_dat_br_lt , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_168 , input \Core_2stage.DatPath_2stage._T , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_1 , input \AsyncScratchPadMemory_2stage.mem_1_MPORT_en , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_ungated_clock , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_15 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_0 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_614 , input \Core_2stage.CtlPath_2stage._csignals_T_99 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_362 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_371 , input \Core_2stage.CtlPath_2stage._csignals_T_57 , input [31:0] io_reset_vector , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_0 , input [31:0] \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_data , input \Core_2stage.DatPath_2stage.csr_io_interrupts_mtip , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_164 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_52 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_7 , input [15:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_7 , input \Core_2stage.d_io_dat_inst_misaligned , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_8 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_225 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_14 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sie , input \Core_2stage.d_io_dat_mem_store , input io_master_port_1_req_valid , input \Core_2stage.DatPath_2stage.csr_io_interrupt , input io_interrupt_meip , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_340 , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_0 , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.value , input \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_0 , input \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_en , input [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_1 , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_1 , input \Core_2stage.CtlPath_2stage.cs0_1 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mie , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugBreak_T_3 , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_1 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_332 , input [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_mask , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_3 , input [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_hi , input \Core_2stage.CtlPath_2stage.io_dat_inst_misaligned , input \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_fcn , input \AsyncScratchPadMemory_2stage.mem_3_MPORT_en , input \Core_2stage.CtlPath_2stage._csignals_T_69 , input [2:0] \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_2 , input [31:0] \AsyncScratchPadMemory_2stage.io_imem_resp_bits_data_state_invariant , input \Core_2stage.DatPath_2stage.CSRFile_2stage._T_222 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_20 , input \Core_2stage.c_io_dat_data_misaligned , input \Core_2stage.DatPath_2stage.csr_io_status_spie , input [31:0] router_1_io_corePort_req_bits_data , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mpie , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_113 , input [31:0] memory_io_core_ports_0_req_bits_data , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_124 , input [31:0] router_1_io_masterPort_req_bits_addr , input \Core_2stage.CtlPath_2stage._csignals_T_37 , input \Core_2stage.CtlPath_2stage._csignals_T_411 , input \Core_2stage.DatPath_2stage.io_ctl_if_kill , input \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_mask , input [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_2 , input [31:0] \Core_2stage.d_io_dat_inst , input [6:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_1 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_599 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_167 , input \Core_2stage.DatPath_2stage.csr_io_csr_stall , input [9:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_addr , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_1 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_3 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_278 , input [62:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._GEN_0 , input router_io_masterPort_resp_valid , input [1:0] \Core_2stage.DatPath_2stage.io_ctl_wb_sel , input \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_en , input [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_3 , input [2:0] \Core_2stage.DatPath_2stage.csr_io_rw_cmd , input [31:0] \Core_2stage.CtlPath_2stage._csignals_T_32 , input [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_vs , input [31:0] \Core_2stage.DatPath_2stage._csr_io_tval_T_6 , input [11:0] \Core_2stage.DatPath_2stage.imm_s , input [31:0] io_master_port_0_req_bits_data , input [32:0] \SodorRequestRouter_2stage_1._in_range_T_3 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_op1_T_4 , input io_master_port_1_resp_valid , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_320 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_28 , input [31:0] \SodorRequestRouter_2stage_0.io_corePort_resp_bits_data , input [31:0] \Core_2stage.DatPath_2stage._if_pc_next_T_5 , input memory_io_core_ports_1_req_valid , input router_io_corePort_resp_valid , input [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_17 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_2 , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_2 , input \Core_2stage.CtlPath_2stage._csignals_T_21 , input \Core_2stage.DatPath_2stage.CSRFile_2stage._T_174 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_269 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_1 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_282 , input [31:0] router_io_masterPort_req_bits_addr , input [31:0] \Core_2stage.DatPath_2stage._tval_inst_ma_T_4 , input [7:0] \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_data , input \Core_2stage.d_io_dat_if_valid_resp , input io_master_port_0_req_bits_fcn , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_636 , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_214 , input [31:0] \Core_2stage.DatPath_2stage.exe_br_target , input [1:0] \Core_2stage.d_io_ctl_mem_fcn , input [9:0] \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_addr , input \Core_2stage.DatPath_2stage._if_pc_next_T_2 , input [31:0] \Core_2stage.DatPath_2stage.exe_alu_out , input \Core_2stage.CtlPath_2stage._csignals_T_13 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_0 , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_maskWithOffset , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_100 , input [31:0] \Core_2stage.DatPath_2stage._csr_io_tval_T_4 , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._sign_T_1 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_237 , input [2:0] \AsyncScratchPadMemory_2stage._io_core_ports_1_resp_bits_data_T_1_state_invariant , input [31:0] \Core_2stage.io_imem_resp_bits_data , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_604 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_19 , input [31:0] \Core_2stage.DatPath_2stage._tval_inst_ma_T_3 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.wdata , input \Core_2stage.CtlPath_2stage._csignals_T_29 , input \Core_2stage.DatPath_2stage.csr_io_status_cease , input router_io_corePort_req_valid , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_wfi , input [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._masks_maskWithOffset_T , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtval , input \Core_2stage.CtlPath_2stage._csignals_T_47 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_606 , input \Core_2stage.DatPath_2stage.csr_io_hartid , input [2:0] \Core_2stage.c_io_ctl_csr_cmd , input [31:0] \Core_2stage.DatPath_2stage._exe_wbdata_T_5 , input \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugTrigger_T_1 , input [2:0] router_io_corePort_req_bits_typ , input [31:0] \Core_2stage.DatPath_2stage._exe_wbdata_T_6 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_107 , input [2:0] \SodorRequestRouter_2stage_0.io_corePort_req_bits_typ , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_108 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_26 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_377 , input [2:0] router_1_io_corePort_req_bits_typ , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.s_offset , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_379 , input [7:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_zero1 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_call , input [1:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_size , input \Core_2stage.DatPath_2stage.csr_io_ungated_clock , input [2:0] \Core_2stage.CtlPath_2stage.io_ctl_pc_sel_no_xept , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus , input [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_fs , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_319 , input [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_1 , input [7:0] \AsyncScratchPadMemory_2stage.mem_3_MPORT_data , input \Core_2stage.CtlPath_2stage.io_dat_mem_store , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_1 , input [10:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_mask_T , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_28 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_1 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_626 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_631 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_108 , input [31:0] \Core_2stage.CtlPath_2stage.io_dat_inst , input \Core_2stage.DatPath_2stage.csr_io_status_wfi , input \Core_2stage.DatPath_2stage._GEN_1 , input router_1_io_corePort_resp_valid , input [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_1 , input [31:0] \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_data , input [30:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_4 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_wdata , input \Core_2stage.CtlPath_2stage.io_dat_br_eq , input \Core_2stage.DatPath_2stage._exe_alu_out_T_16 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_120 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._m_interrupts_T_3 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_op2_T_5 , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_219 , input [31:0] \Core_2stage.DatPath_2stage.regfile_5 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_210 , input [9:0] \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_addr , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_105 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sd_rv32 , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_1 , input [2:0] \Core_2stage.d_io_ctl_csr_cmd , input [2:0] \Core_2stage.c_io_ctl_pc_sel_no_xept , input [9:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_addr , input \Core_2stage.DatPath_2stage.CSRFile_2stage._T_14 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.system_insn , input \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_0 , input \Core_2stage.CtlPath_2stage._csignals_T_537 , input [6:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_0 , input \Core_2stage.CtlPath_2stage.stall , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_118 , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_114 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_125 , input [31:0] \Core_2stage.DatPath_2stage.regfile_8 , input \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_215 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_197 , input \Core_2stage.DatPath_2stage.regfile_MPORT_mask , input [31:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_data , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_191 , input \Core_2stage.DatPath_2stage.csr_io_status_mprv , input [31:0] \Core_2stage.DatPath_2stage.regfile_12 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_224 , input \Core_2stage.DatPath_2stage._exe_alu_op2_T_2 , input [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_3 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_33 , input \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_fcn , input memory_io_core_ports_0_req_valid , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_23 , input [7:0] \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_data , input [1:0] \Core_2stage.c_io_ctl_wb_sel , input \Core_2stage.CtlPath_2stage._csignals_T_73 , input \AsyncScratchPadMemory_2stage.mem_3_MPORT_mask , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_1 , input [31:0] \SodorRequestRouter_2stage_1.io_masterPort_resp_bits_data , input \Core_2stage.CtlPath_2stage._csignals_T_43 , input [62:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._shiftedVec_T_1 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_21 , input [2:0] \SodorRequestRouter_2stage_1.io_masterPort_req_bits_typ , input [20:0] \AsyncScratchPadMemory_2stage.module__io_addr , input \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_3 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_18 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_239 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_12 , input \Core_2stage.CtlPath_2stage._csignals_T_65 , input [4:0] \Core_2stage.DatPath_2stage.exe_rs1_addr , input \Core_2stage.CtlPath_2stage.io_ctl_mem_val , input \Core_2stage.io_hartid , input [31:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_18 , input \AsyncScratchPadMemory_2stage.mem_2_MPORT_mask , input \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_en , input \Core_2stage.CtlPath_2stage.cs0_0 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_589 , input \Core_2stage.DatPath_2stage._T_1 , input [31:0] \Core_2stage.DatPath_2stage.regfile_27 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_344 , input \Core_2stage.d_io_ctl_exception , input [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_5 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_598 , input [31:0] \Core_2stage.io_reset_vector , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_342 , input [11:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.debugTVec , input \Core_2stage.DatPath_2stage._exe_alu_out_T_17 , input \Core_2stage.DatPath_2stage.CSRFile_2stage._T_367 , input [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_11 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_cease , input [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_0 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_step , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_207 , input router_io_masterPort_req_valid , input [6:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._GEN_1 , input \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_3 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_2 , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._bytes_T_3 , input [3:0] \Core_2stage.CtlPath_2stage.cs_br_type , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_244 , input [9:0] \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_addr , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_19 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_gva , input \Core_2stage.CtlPath_2stage._csignals_T_9 , input \Core_2stage.CtlPath_2stage._csignals_T_130 , input \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_fcn , input \Core_2stage.DatPath_2stage.io_dat_br_eq , input \AsyncScratchPadMemory_2stage.module__io_mem_masks_0 , input io_master_port_0_resp_valid , input \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_51 , input \Core_2stage.DatPath_2stage.csr_io_status_gva , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_205 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_381 , input [2:0] \SodorRequestRouter_2stage_0.io_masterPort_req_bits_typ , input \Core_2stage.DatPath_2stage.io_ctl_stall , input [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._masks_maskWithOffset_T , input [31:0] \Core_2stage.DatPath_2stage.tval_inst_ma , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_ube , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_112 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_2 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_273 , input [1:0] \Core_2stage.DatPath_2stage.csr_io_status_uxl , input \Core_2stage.DatPath_2stage.csr_io_status_sd_rv32 , input [31:0] \Core_2stage.io_imem_req_bits_addr_state_invariant , input [31:0] \Core_2stage.DatPath_2stage.io_imem_resp_bits_data_state_invariant , input \Core_2stage.CtlPath_2stage.io_dmem_req_valid , input \Core_2stage.CtlPath_2stage._csignals_T_540 , input [31:0] \Core_2stage.DatPath_2stage.regfile_30 , input [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_218 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dscratch , input memory_io_debug_port_resp_valid , input [7:0] \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_data , input [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T , input \Core_2stage.d_io_imem_resp_valid , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_108 , input [6:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.nextSmall_1 , input [2:0] memory_io_core_ports_0_req_bits_typ , input \Core_2stage.CtlPath_2stage._csignals_T_67 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_609 , input \Core_2stage.DatPath_2stage.CSRFile_2stage._T_186 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_633 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_cause , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_3 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._cause_T_5 , input \SodorRequestRouter_2stage_1.io_corePort_req_valid , input memory_clock , input \AsyncScratchPadMemory_2stage.mem_0_MPORT_en , input \Core_2stage.DatPath_2stage.csr_io_status_hie , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_1 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_369 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_211 , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_218 , input [1:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_size , input \Core_2stage.CtlPath_2stage._csignals_T_45 , input [1:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_size_state_invariant , input [31:0] \Core_2stage.io_dmem_req_bits_data , input router_io_scratchPort_req_valid , input \Core_2stage.CtlPath_2stage._csignals_T_539 , input [31:0] \Core_2stage.DatPath_2stage.regfile_21 , input [31:0] \Core_2stage.DatPath_2stage.exe_reg_pc , input \Core_2stage.CtlPath_2stage.io_dat_csr_eret , input \Core_2stage.DatPath_2stage.csr_clock , input [31:0] \SodorRequestRouter_2stage_1.io_masterPort_req_bits_addr , input [31:0] \Core_2stage.CtlPath_2stage._csignals_T_16 , input \Core_2stage.DatPath_2stage.CSRFile_2stage._io_interrupt_T , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_18 , input [4:0] \Core_2stage.DatPath_2stage.io_ctl_alu_fun , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_128 , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_1 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_277 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_40 , input [19:0] \Core_2stage.DatPath_2stage._imm_s_sext_T_2 , input \Core_2stage.DatPath_2stage._GEN_3 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_28 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_1 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.csr_wen , input \SodorRequestRouter_2stage_1.io_scratchPort_resp_valid , input [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_1 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_36 , input \Core_2stage.DatPath_2stage._if_pc_next_T , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_38 , input core_io_hartid , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sbe , input [31:0] \Core_2stage.DatPath_2stage.io_dmem_req_bits_addr , input [2:0] io_master_port_0_req_bits_typ , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_15 , input \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_2 , input \Core_2stage.DatPath_2stage.io_dat_br_lt , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_12 , input [31:0] router_1_io_scratchPort_req_bits_data , input [31:0] \Core_2stage.DatPath_2stage.regfile_0 , input [2:0] \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_typ , input \Core_2stage.CtlPath_2stage.io_dat_if_valid_resp , input [31:0] \SodorRequestRouter_2stage_0.io_corePort_req_bits_data , input \Core_2stage.CtlPath_2stage._csignals_T_7 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_2 , input [1:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_size , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_singleStepped , input [4:0] \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_addr , input [31:0] io_master_port_1_req_bits_addr , input [31:0] \Core_2stage.d_io_imem_resp_bits_data , input [31:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_data , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_2 , input [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_2_state_invariant , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_98 , input [1:0] \Core_2stage.DatPath_2stage.csr_io_status_xs , input \Core_2stage.CtlPath_2stage._csignals_T_41 , input [4:0] \Core_2stage.DatPath_2stage.exe_wbaddr , input \SodorRequestRouter_2stage_1.resp_in_range , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_115 , input [7:0] \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_data , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_41 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_170 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_338 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease_r , input [31:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_req_bits_addr , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_310 , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.bytes , input [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_2 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_211 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_279 , input [31:0] \Core_2stage.DatPath_2stage.regfile_31 , input [2:0] \Core_2stage.d_io_ctl_pc_sel_no_xept , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_387 , input [1:0] \Core_2stage.DatPath_2stage.csr_io_status_prv , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_304 , input \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_valid , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_352 , input [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcountinhibit , input \Core_2stage.c_io_dmem_req_valid , input \Core_2stage.DatPath_2stage._exe_alu_op1_T_1 , input [7:0] \AsyncScratchPadMemory_2stage.module__io_mem_data_2 , input \Core_2stage.io_imem_req_valid , input [2:0] \Core_2stage.CtlPath_2stage.io_ctl_op2_sel , input \Core_2stage.d_reset , input \Core_2stage.DatPath_2stage.io_dat_if_valid_resp , input [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._masks_maskWithOffset_T , input \Core_2stage.CtlPath_2stage.cs_val_inst , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_10 , input [20:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_addr , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_2 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_3 , input [31:0] \Core_2stage.DatPath_2stage.io_imem_resp_bits_data , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_34 , input \Core_2stage.CtlPath_2stage._csignals_T_407 , input [31:0] \Core_2stage.DatPath_2stage.exe_rs2_data , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_2 , input [9:0] \AsyncScratchPadMemory_2stage.mem_0_MPORT_addr , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_size , input [5:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_35 , input \Core_2stage.CtlPath_2stage.io_dat_br_ltu , input [31:0] router_io_scratchPort_req_bits_data , input [31:0] \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_addr , input [31:0] \Core_2stage.DatPath_2stage.regfile_20 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_174 , input [10:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_mask_T , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_18 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mepc , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_1 , input \Core_2stage.d_clock , input \Core_2stage.DatPath_2stage._csr_io_tval_T_1 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_603 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec , input [31:0] \Core_2stage.DatPath_2stage.if_pc_plus4 , input \SodorRequestRouter_2stage_1.in_range , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_182 , input [31:0] \Core_2stage.DatPath_2stage._io_dat_br_lt_T_1 , input \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_fcn , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_97 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_318 , input [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_2 , input \Core_2stage.CtlPath_2stage._csignals_T_19 , input [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_1 , input [3:0] \Core_2stage.CtlPath_2stage.cs_alu_fun , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_267 , input \Core_2stage.CtlPath_2stage._csignals_T_53 , input [1:0] \Core_2stage.DatPath_2stage.io_ctl_mem_fcn , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_3 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_271 , input \Core_2stage.io_dmem_resp_valid , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.m_interrupts , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_csr_stall , input \Core_2stage.CtlPath_2stage._csignals_T_15 , input [31:0] \Core_2stage.DatPath_2stage.regfile_MPORT_1_data , input \Core_2stage.DatPath_2stage.csr_reset , input \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_242 , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_120 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_333 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_634 , input \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_en , input [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_3 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_1 , input [31:0] io_master_port_1_req_bits_data , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_31 , input [31:0] \SodorRequestRouter_2stage_1._in_range_T , input [31:0] \Core_2stage.DatPath_2stage.imm_j_sext , input \Core_2stage.c_io_dat_inst_misaligned , input \Core_2stage.DatPath_2stage.csr_io_status_debug , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_179 , input [2:0] \Core_2stage.CtlPath_2stage.io_ctl_pc_sel , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_6 , input \Core_2stage.CtlPath_2stage._csignals_T_17 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_228 , input [20:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_addr , input [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_216 , input [2:0] \AsyncScratchPadMemory_2stage._io_core_ports_0_resp_bits_data_T_1 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.epc , input [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_3 , input [2:0] \Core_2stage.DatPath_2stage._io_dat_data_misaligned_T_1 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_334 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_9 , input [5:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.small_1 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_289 , input \SodorRequestRouter_2stage_0.io_corePort_req_bits_fcn , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.s_offset , input memory_io_core_ports_0_resp_valid , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_2 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_12 , input \Core_2stage.DatPath_2stage.reset , input \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_3 , input [2:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_typ , input \Core_2stage.DatPath_2stage.csr_io_status_sd , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_638 , input [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._masks_maskWithOffset_T , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_173 , input \Core_2stage.d_io_ctl_mem_val , input [2:0] router_1_io_masterPort_req_bits_typ , input [31:0] \Core_2stage.DatPath_2stage.regfile_10 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_384 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_uie , input [9:0] \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_addr , input \Core_2stage.DatPath_2stage._exe_alu_out_T_15 , input [9:0] \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_addr , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_0 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_355 , input \Core_2stage.DatPath_2stage.csr_io_status_mpie , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_size , input \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_1 , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_28 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_11 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_175 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_331 , input core_io_dmem_req_valid , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_23 , input core_io_interrupt_debug , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_5 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_pc , input router_1_io_scratchPort_req_valid , input \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_180 , input [9:0] \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_addr , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_time , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.addr , input [31:0] \Core_2stage.DatPath_2stage.regfile_9 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_290 , input [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_maskWithOffset , input [31:0] \SodorRequestRouter_2stage_0.io_corePort_req_bits_addr , input [2:0] \Core_2stage.DatPath_2stage._misaligned_mask_T_1 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_372 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_12 , input \Core_2stage.DatPath_2stage.csr_io_status_mbe , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mprv , input [2:0] \Core_2stage.c_io_ctl_pc_sel , input [2:0] router_1_io_scratchPort_req_bits_typ , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_233 , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.bytes , input [7:0] \AsyncScratchPadMemory_2stage.mem_0_MPORT_data , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo , input [31:0] \Core_2stage.DatPath_2stage.imm_b_sext , input [11:0] \Core_2stage.DatPath_2stage.csr_io_rw_addr , input [2:0] \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T , input \Core_2stage.c_io_ctl_mem_val , input \Core_2stage.io_dmem_req_bits_fcn , input \SodorRequestRouter_2stage_0.io_scratchPort_resp_valid , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1719 , input [9:0] \AsyncScratchPadMemory_2stage.module_1_io_mem_addr , input memory_io_debug_port_req_bits_fcn , input \Core_2stage.reset , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_386 , input [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_2 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_3 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_268 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_595 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_588 , input [31:0] \Core_2stage.DatPath_2stage.pc_x , input [31:0] \Core_2stage.DatPath_2stage._T_4 , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_2 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_op1_T_3 , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._bytes_T_1 , input \Core_2stage.DatPath_2stage.io_imem_resp_valid , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_117 , input [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_2 , input [2:0] \Core_2stage.DatPath_2stage.io_ctl_pc_sel , input \SodorRequestRouter_2stage_0.io_masterPort_resp_valid , input \Core_2stage.DatPath_2stage.csr_io_status_dv , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_315 , input \Core_2stage.DatPath_2stage.io_interrupt_mtip , input [32:0] \SodorRequestRouter_2stage_0._in_range_T_1 , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._bytes_T_3 , input [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_207 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_4 , input [7:0] \AsyncScratchPadMemory_2stage.module_1_io_mem_data_3 , input \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_3 , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_118 , input [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_0_state_invariant , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_630 , input \Core_2stage.CtlPath_2stage._csignals_T_438 , input \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_signed , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_7 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_2 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_2 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_1 , input [9:0] \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_addr , input \Core_2stage.d_io_dat_csr_interrupt , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_2 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_31 , input \Core_2stage.CtlPath_2stage.io_ctl_rf_wen , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_2 , input [1:0] \Core_2stage.CtlPath_2stage.io_ctl_mem_fcn , input [31:0] \SodorRequestRouter_2stage_0.io_masterPort_resp_bits_data , input \Core_2stage.DatPath_2stage.io_interrupt_msip , input [31:0] \Core_2stage.DatPath_2stage.regfile_22 , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_103 , input \Core_2stage.DatPath_2stage._exe_alu_out_T_6 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_173 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_374 , input [31:0] \Core_2stage.DatPath_2stage.exe_alu_op1 , input \Core_2stage.CtlPath_2stage._csignals_T_83 , input [31:0] \Core_2stage.DatPath_2stage._exe_jump_reg_target_T_1 , input \AsyncScratchPadMemory_2stage.module_1_io_en , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.bytes , input \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_241 , input [2:0] \Core_2stage.c_io_ctl_op2_sel , input [64:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_hi_hi , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_341 , input \Core_2stage.DatPath_2stage._exe_wbdata_T , input \Core_2stage.CtlPath_2stage.io_dat_br_lt , input \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_279 , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._bytes_T_3 , input \SodorRequestRouter_2stage_1.io_corePort_resp_valid , input \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_signed , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_2 , input [31:0] \Core_2stage.DatPath_2stage.csr_io_status_isa , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_194 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpv , input \Core_2stage.DatPath_2stage._csr_io_tval_T , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_102 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_325 , input \Core_2stage.DatPath_2stage.exe_wben , input \Core_2stage.DatPath_2stage.io_ctl_rf_wen , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_287 , input [31:0] \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_data , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_628 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_10 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_176 , input [31:0] \Core_2stage.DatPath_2stage.regfile_26 , input [31:0] \Core_2stage.CtlPath_2stage.io_ctl_exception_cause , input [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_2 , input [31:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_data , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_27 , input memory_io_core_ports_0_req_bits_fcn , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_209 , input [31:0] \Core_2stage.DatPath_2stage.exe_jump_reg_target , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_size , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_585 , input [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_0 , input [31:0] \Core_2stage.DatPath_2stage.regfile_24 , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.whichInterrupt , input [31:0] \Core_2stage.DatPath_2stage.regfile_29 , input \Core_2stage.DatPath_2stage._exe_alu_out_T_18 , input \Core_2stage.CtlPath_2stage.io_dmem_req_bits_fcn , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_232 , input [4:0] \Core_2stage.d_io_ctl_alu_fun , input \Core_2stage.DatPath_2stage.CSRFile_2stage._T_180 , input [7:0] \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_data , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_356 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_600 , input [31:0] \Core_2stage.DatPath_2stage.regfile_6 , input [4:0] \Core_2stage.CtlPath_2stage.rs1_addr , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_107 , input [4:0] \Core_2stage.DatPath_2stage.regfile_MPORT_1_addr , input [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_lo , input [31:0] \Core_2stage.DatPath_2stage.regfile_17 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tvm , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_11 , input \Core_2stage.DatPath_2stage.csr_io_status_mie , input [31:0] \SodorRequestRouter_2stage_1.io_corePort_req_bits_addr , input [20:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_addr , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_234 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T , input [31:0] \Core_2stage.DatPath_2stage.imm_u_sext , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_28 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_4 , input router_io_corePort_req_bits_fcn , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_op2_T_4 , input [9:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_addr , input [31:0] \Core_2stage.DatPath_2stage.csr_io_time , input [31:0] \Core_2stage.DatPath_2stage._if_pc_next_T_7 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_162 , input \Core_2stage.DatPath_2stage.csr_io_singleStep , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_388 , input [31:0] memory_io_debug_port_resp_bits_data , input \Core_2stage.DatPath_2stage.CSRFile_2stage.anyInterrupt , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_32 , input [31:0] \Core_2stage.DatPath_2stage.csr_io_tval , input [31:0] \Core_2stage.DatPath_2stage.csr_io_rw_wdata , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_357 , input memory_io_debug_port_req_valid , input [31:0] memory_io_core_ports_0_req_bits_addr , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_1 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_241 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease , input \Core_2stage.DatPath_2stage.CSRFile_2stage.exception , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_122 , input \Core_2stage.DatPath_2stage.regfile_MPORT_en , input [31:0] \AsyncScratchPadMemory_2stage.module_1_io_data , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_339 , input [31:0] \SodorRequestRouter_2stage_0._resp_in_range_T , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_337 , input [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_23 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_4 , input \Core_2stage.DatPath_2stage.clock , input [31:0] \Core_2stage.DatPath_2stage.regfile_28 , input [2:0] \Core_2stage.c_io_dmem_req_bits_typ , input \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_en , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_190 , input [1:0] \Core_2stage.c_io_ctl_mem_fcn , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_235 , input \Core_2stage.DatPath_2stage._exe_alu_out_T_3 , input [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_1 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_635 , input [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_lo , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_2 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_20 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sd , input [31:0] router_io_corePort_req_bits_addr , input [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_293 , input \Core_2stage.DatPath_2stage._if_pc_next_T_1 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_27 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_28 , input \Core_2stage.DatPath_2stage.csr_io_status_spp , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_14 , input [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sxl , input [32:0] \SodorRequestRouter_2stage_0._resp_in_range_T_3 , input [7:0] \AsyncScratchPadMemory_2stage.module__io_mem_data_1 , input \Core_2stage.DatPath_2stage._exe_alu_op2_T , input [19:0] \Core_2stage.DatPath_2stage.imm_u , input [2:0] \AsyncScratchPadMemory_2stage._io_debug_port_resp_bits_data_T_1 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_0 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_389 , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_300 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_1 , input [31:0] \SodorRequestRouter_2stage_0.io_respAddress , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_323 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_620 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_0 , input [31:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_data , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_283 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mie , input \Core_2stage.DatPath_2stage.if_inst_buffer_valid , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_2 , input \Core_2stage.CtlPath_2stage._csignals_T_409 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_593 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_584 , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_104 , input [1:0] \Core_2stage.DatPath_2stage.io_ctl_op1_sel , input \Core_2stage.DatPath_2stage.io_interrupt_meip , input \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_en , input [7:0] \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_data , input [14:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.d_interrupts , input [31:0] router_io_scratchPort_resp_bits_data , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_36 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_188 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_632 , input [1:0] \Core_2stage.CtlPath_2stage.io_ctl_op1_sel , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_116 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_329 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_216 , input router_io_scratchPort_req_bits_fcn , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_2 , input core_io_interrupt_msip , input [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_3_state_invariant , input \Core_2stage.DatPath_2stage.csr_io_status_ube , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_183 , input \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugInt_T_1 , input \Core_2stage.DatPath_2stage.csr_io_status_sie , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_177 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_doVector , input [2:0] memory_io_debug_port_req_bits_typ , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._bytes_T_1 , input \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.sign , input [6:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.nextSmall , input \Core_2stage.DatPath_2stage.io_interrupt_debug , input [20:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_addr , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_12 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_213 , input [31:0] \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_data , input \Core_2stage.CtlPath_2stage._csignals_T_3 , input \Core_2stage.CtlPath_2stage._csignals_T_39 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mie_T , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_19 , input [31:0] \Core_2stage.DatPath_2stage.csr_io_evec , input [2:0] \Core_2stage.CtlPath_2stage.ctrl_pc_sel , input [7:0] \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_data , input \Core_2stage.DatPath_2stage.io_ctl_exception , input [1:0] \Core_2stage.DatPath_2stage.csr_io_status_vs , input [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_13 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_305 , input [31:0] \Core_2stage.DatPath_2stage.io_imem_req_bits_addr , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._m_interrupts_T_5 , input [32:0] \SodorRequestRouter_2stage_0._resp_in_range_T_1 , input [31:0] \Core_2stage.DatPath_2stage.imm_i_sext , input [31:0] io_debug_port_req_bits_data , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_3 , input [31:0] \Core_2stage.DatPath_2stage.regfile_13 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_1 , input [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpp , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_evec , input \Core_2stage.DatPath_2stage.CSRFile_2stage._T_366 , input [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_1 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_239 , input [31:0] memory_io_debug_port_req_bits_addr , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_623 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_0 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_608 , input \Core_2stage.DatPath_2stage.csr_io_interrupts_meip , input \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_1 , input \Core_2stage.DatPath_2stage.decode , input [31:0] \Core_2stage.DatPath_2stage.exe_reg_inst , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_318 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_124 , input io_debug_port_req_bits_fcn , input [31:0] \AsyncScratchPadMemory_2stage.io_imem_req_bits_addr_state_invariant , input [31:0] \Core_2stage.DatPath_2stage.exe_alu_op2 , input [2:0] router_io_scratchPort_req_bits_typ , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_303 , input [31:0] memory_io_debug_port_req_bits_data , input \AsyncScratchPadMemory_2stage.io_core_ports_1_req_valid , input \Core_2stage.DatPath_2stage.io_hartid , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_341 , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_18 , input \Core_2stage.DatPath_2stage.csr_io_status_tw , input [9:0] \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_addr , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1717 , input [2:0] \Core_2stage.DatPath_2stage.misaligned_mask , input [32:0] \SodorRequestRouter_2stage_0._in_range_T_3 , input \Core_2stage.CtlPath_2stage.csr_ren , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_213 , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_129 , input [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_1 , input [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_26 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_11 , input io_interrupt_debug , input [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T , input \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_48 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_172 , input [62:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._shiftedVec_T_1 , input [31:0] \Core_2stage.DatPath_2stage._io_dat_br_lt_T , input [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_22 , input \Core_2stage.CtlPath_2stage.illegal , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_296 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_218 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_613 , input \Core_2stage.c_io_dat_br_lt , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_317 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_354 , input [31:0] core_io_dmem_req_bits_addr , input [31:0] \SodorRequestRouter_2stage_1._resp_in_range_T , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.bytes , input [7:0] \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_data , input \Core_2stage.CtlPath_2stage._csignals_T_35 , input \Core_2stage.DatPath_2stage.csr_io_status_mxr , input \Core_2stage.CtlPath_2stage._csignals_T_75 , input [5:0] \Core_2stage.DatPath_2stage._misaligned_mask_T_4 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_7 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_169 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_326 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_3 , input [7:0] \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_data , input router_1_io_scratchPort_resp_valid , input \Core_2stage.CtlPath_2stage._csignals_T_59 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_605 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_0 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_rdata , input [31:0] \Core_2stage.io_dmem_req_bits_addr , input \Core_2stage.CtlPath_2stage._csignals_T_23 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcause , input io_debug_port_resp_valid , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_12 , input \Core_2stage.clock , input [2:0] \Core_2stage.DatPath_2stage.io_ctl_op2_sel , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_166 , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_130 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_174 , input [31:0] \Core_2stage.DatPath_2stage.imm_s_sext , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_242 , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.cause , input [31:0] \Core_2stage.DatPath_2stage.exe_rs1_data , input \Core_2stage.CtlPath_2stage._csignals_T_25 , input [1:0] \AsyncScratchPadMemory_2stage.module_1_io_size , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_360 , input [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_20 , input [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_1 , input [7:0] \AsyncScratchPadMemory_2stage.module__io_mem_data_3 , input \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_en , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_19 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_594 , input [19:0] \Core_2stage.DatPath_2stage.imm_j , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_270 , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._sign_T_1 , input io_debug_port_req_valid , input [31:0] io_imem_resp_bits_data_state_invariant , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_212 , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1714 , input \Core_2stage.io_dmem_req_valid , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_22 , input [4:0] \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_addr , input [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T , input \AsyncScratchPadMemory_2stage.mem_0_MPORT_mask , input [31:0] \Core_2stage.DatPath_2stage.io_imem_req_bits_addr_state_invariant , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_176 , input [9:0] \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_addr , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_272 , input [31:0] \Core_2stage.c_io_dat_inst , input [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_18 , input \Core_2stage.DatPath_2stage.csr_io_interrupts_msip , input [1:0] \AsyncScratchPadMemory_2stage.module__io_size , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_336 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_2 , input \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_2 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_186 , input [31:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_96 , input core_reset , input \AsyncScratchPadMemory_2stage.io_core_ports_0_req_valid , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_343 , input [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_18 , input [31:0] \Core_2stage.DatPath_2stage._csr_io_tval_T_5 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_308 , input \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_6 , input [31:0] \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_data , input [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_0 , input [31:0] \Core_2stage.d_io_dmem_req_bits_addr , input \Core_2stage.DatPath_2stage.CSRFile_2stage._T_177 , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_629 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_311 , input [6:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_maskWithOffset_T , input [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_lo , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_230 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_16 , input [1:0] \Core_2stage.DatPath_2stage.csr_io_status_dprv , input [31:0] \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_addr , input [7:0] \AsyncScratchPadMemory_2stage.module__io_mem_data_0 , input [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_24 , input [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_xs , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_7 , input \Core_2stage.c_io_ctl_if_kill , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_3 , input [9:0] \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_addr , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_1 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_163 , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_597 , input [31:0] \Core_2stage.DatPath_2stage.regfile_16 , input core_io_dmem_resp_valid , input \Core_2stage.DatPath_2stage.io_dat_csr_interrupt , input \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_signed , input \SodorRequestRouter_2stage_1.io_masterPort_req_valid , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_182 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_366 , input [31:0] core_io_imem_resp_bits_data , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_10 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_19 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_165 , input \Core_2stage.io_interrupt_debug , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_4 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_0 , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_375 , input [31:0] \SodorRequestRouter_2stage_0._in_range_T , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_1 , input \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_en , input \Core_2stage.DatPath_2stage.CSRFile_2stage.x79 , input [2:0] \Core_2stage.CtlPath_2stage.io_ctl_csr_cmd , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_5 , input \Core_2stage.io_imem_resp_valid , input [7:0] \Core_2stage.DatPath_2stage._T_14 , input io_hartid , input [1:0] \Core_2stage.d_io_ctl_wb_sel , input [31:0] \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_addr , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_382 , input [20:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_addr , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_eret , input \Core_2stage.DatPath_2stage.csr_io_status_tsr , input [11:0] \Core_2stage.DatPath_2stage.imm_i , input [31:0] \Core_2stage.CtlPath_2stage._csignals_T , input [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_122 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_185 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_6 , input [11:0] \Core_2stage.DatPath_2stage.imm_b , input [2:0] \Core_2stage.DatPath_2stage.io_ctl_mem_typ , input \Core_2stage.DatPath_2stage.regfile_MPORT_1_en , input \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_en , input \Core_2stage.DatPath_2stage.io_dat_inst_misaligned , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_612 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_171 , input \Core_2stage.CtlPath_2stage._csignals_T_89 , input \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_46 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_spp , input [2:0] \Core_2stage.CtlPath_2stage._csignals_T_288 , input [1:0] \Core_2stage.CtlPath_2stage.io_ctl_wb_sel , input [31:0] router_1_io_respAddress , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_214 , input \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_en , input [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_2 , input router_io_scratchPort_resp_valid , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reset , input \SodorRequestRouter_2stage_1.io_masterPort_resp_valid , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_9 , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_v , input [1:0] \Core_2stage.CtlPath_2stage._csignals_T_391 , input [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_95 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_180 , input \Core_2stage.CtlPath_2stage.io_ctl_if_kill , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_314 , input [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_298 , input \Core_2stage.CtlPath_2stage._csignals_T_412 , input [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_20 , input \Core_2stage.DatPath_2stage.exe_reg_valid , input [7:0] \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_data , input [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._sign_T_1 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_189 , input [3:0] \Core_2stage.CtlPath_2stage._csignals_T_330 , input \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_en , input \Core_2stage.DatPath_2stage._exe_alu_out_T_10 , input [31:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_addr , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_7_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_reset_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_data_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_216_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_16_obs_trg_cond , output \Core_2stage.DatPath_2stage._imm_s_sext_T_2_obs_trg_cond , output \Core_2stage.c_io_ctl_if_kill_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_19_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.epc_obs_trg_arg0 , output \Core_2stage.c_io_ctl_mem_typ_obs_trg_cond , output \Core_2stage.DatPath_2stage._csr_io_tval_T_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_38_obs_trg_cond , output router_io_scratchPort_req_valid_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_114_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.cause_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_cease_obs_trg_cond , output [31:0] \SodorRequestRouter_2stage_1.io_masterPort_req_bits_addr_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_619_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_0_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_107_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_34_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_614_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_106_obs_trg_cond , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_18_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_17_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_122_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_1_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_292_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_fcn_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._if_pc_next_T_5_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_6_obs_trg_cond , output [1:0] \Core_2stage.DatPath_2stage.csr_io_status_fs_obs_trg_arg0 , output \Core_2stage.d_io_imem_req_bits_addr_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_spie_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.module_1_io_mem_data_2_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_325_obs_trg_cond , output router_1_io_masterPort_req_bits_fcn_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_vs_obs_trg_arg0 , output \Core_2stage.d_io_interrupt_msip_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_exception_obs_trg_cond , output [20:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_addr_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_2_obs_trg_cond , output [31:0] io_master_port_0_req_bits_addr_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_266_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_32_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_uxl_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_34_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_exception_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_178_obs_trg_cond , output [31:0] io_debug_port_req_bits_addr_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.module__io_en_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._masks_maskWithOffset_T_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_11_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_ctl_csr_cmd_obs_trg_cond , output [31:0] \SodorRequestRouter_2stage_0.io_masterPort_req_bits_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.new_mstatus_mpie_obs_trg_cond , output \SodorRequestRouter_2stage_1.io_masterPort_req_bits_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_debug_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_27_obs_trg_cond , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_268_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_mtip_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.s_offset_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_debug_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_1_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_315_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_213_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_1_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_126_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_tval_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_615_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_doVector_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.bytes_obs_trg_arg0 , output io_master_port_1_resp_valid_obs_trg_cond , output \SodorRequestRouter_2stage_1.resp_in_range_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_5_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_8_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.exe_alu_op1_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_arg0 , output [18:0] \Core_2stage.DatPath_2stage._imm_b_sext_T_2_obs_trg_arg0 , output [31:0] core_io_dmem_req_bits_addr_obs_trg_arg0 , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_obs_trg_arg0 , output memory_io_debug_port_req_bits_fcn_obs_trg_cond , output \SodorRequestRouter_2stage_1._resp_in_range_T_3_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.exe_alu_out_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._any_T_78_obs_trg_cond , output [104:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mstatus_T_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_51_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.in_range_obs_trg_cond , output \Core_2stage.c_io_dmem_req_valid_obs_trg_cond , output \Core_2stage.DatPath_2stage._GEN_1_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tw_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_dat_csr_interrupt_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_3_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_en_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_185_obs_trg_arg0 , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_38_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_538_obs_trg_arg0 , output [32:0] \SodorRequestRouter_2stage_0._in_range_T_3_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_hi_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_ube_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_1_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_112_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._exe_wbdata_T_4_obs_trg_arg0 , output [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_maskWithOffset_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_19_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_286_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_size_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_438_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_113_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_27_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_381_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_243_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_hi_hi_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_583_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_121_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_598_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_1_obs_trg_cond , output \SodorRequestRouter_2stage_1.io_corePort_req_bits_fcn_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_9_obs_trg_arg0 , output [2:0] io_master_port_1_req_bits_typ_obs_trg_arg0 , output [31:0] router_1_io_corePort_req_bits_addr_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_274_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_0_obs_trg_cond , output [31:0] router_1_io_masterPort_req_bits_addr_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_378_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_107_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_op2_T_1_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.exe_jump_reg_target_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_upie_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.bytes_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_dat_data_misaligned_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_arg0 , output router_1_io_scratchPort_req_bits_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_593_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_en_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_2_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.rs1_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugBreak_obs_trg_arg0 , output [2:0] \Core_2stage.DatPath_2stage.io_ctl_mem_typ_obs_trg_arg0 , output [2:0] \Core_2stage.c_io_ctl_mem_typ_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_0_obs_trg_cond , output \Core_2stage.DatPath_2stage._GEN_1_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_12_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_114_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_601_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_43_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_size_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_167_obs_trg_cond , output [5:0] \Core_2stage.DatPath_2stage._misaligned_mask_T_3_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1717_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_24_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._large_r_T_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_wfi_obs_trg_cond , output io_master_port_0_req_bits_fcn_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.exe_reg_pc_plus4_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.io_dmem_req_bits_addr_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_3_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_addr_obs_trg_arg0 , output \Core_2stage.c_io_dmem_req_valid_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_382_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_respAddress_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_spie_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_174_obs_trg_arg0 , output INSTR_inv_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_2_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.module__io_mem_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tsr_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_3_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_225_obs_trg_cond , output [4:0] \Core_2stage.DatPath_2stage.regfile_MPORT_1_addr_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.csr_ren_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_335_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_307_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_addr_obs_trg_cond , output \Core_2stage.d_io_ctl_exception_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_3_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_228_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_dat_inst_obs_trg_cond , output [31:0] router_1_io_scratchPort_resp_bits_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_27_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_326_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_31_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_9_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_dmem_resp_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_csr_stall_obs_trg_cond , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_117_obs_trg_arg0 , output [7:0] \Core_2stage.DatPath_2stage._T_17_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_11_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_2_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_384_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_12_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage.io_ctl_pc_sel_no_xept_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_exception_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_upie_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_singleStepped_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_234_obs_trg_arg0 , output router_io_corePort_req_bits_typ_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._shiftedVec_T_obs_trg_cond , output \Core_2stage.io_dmem_req_bits_data_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_128_obs_trg_arg0 , output [31:0] memory_io_core_ports_0_resp_bits_data_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.whichInterrupt_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_30_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_26_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_retire_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_masterPort_req_bits_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.exe_reg_inst_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_27_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_52_obs_trg_arg0 , output \Core_2stage.io_interrupt_msip_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_337_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_2_obs_trg_cond , output [2:0] \Core_2stage.d_io_ctl_mem_typ_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_187_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_30_obs_trg_cond , output [31:0] memory_io_debug_port_req_bits_data_obs_trg_arg0 , output [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_lo_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_data_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.module__io_mem_masks_0_obs_trg_arg0 , output [31:0] core_io_dmem_resp_bits_data_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_3_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_dat_br_eq_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_176_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_333_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_break_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_16_obs_trg_arg0 , output [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_maskWithOffset_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_data_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_228_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_break_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_237_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_1_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.tval_inst_ma_obs_trg_arg0 , output \Core_2stage.d_io_dat_br_lt_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_pc_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_10_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._any_T_78_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_116_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_interrupts_msip_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_22_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mie_obs_trg_cond , output [2:0] \AsyncScratchPadMemory_2stage._io_debug_port_resp_bits_data_T_1_obs_trg_arg0 , output [30:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_4_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_masterPort_req_bits_addr_obs_trg_cond , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_22_obs_trg_arg0 , output [20:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_addr_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_173_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._if_pc_next_T_7_obs_trg_arg0 , output RDATA_inv_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_341_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module__io_mem_data_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mscratch_obs_trg_cond , output \SodorRequestRouter_2stage_0._resp_in_range_T_3_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_data_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_2_obs_trg_arg0 , output \Core_2stage.c_io_dmem_req_bits_typ_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_1_obs_trg_cond , output [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_59_obs_trg_arg0 , output [31:0] router_io_corePort_req_bits_addr_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_2_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_28_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_hie_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mbe_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_obs_trg_cond , output [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_maskWithOffset_obs_trg_arg0 , output router_1_io_masterPort_resp_bits_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_1_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.new_mstatus_mpie_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.mem_2_MPORT_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_97_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_146_obs_trg_cond , output \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_2_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_236_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_31_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_222_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_size_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage.io_ctl_op2_sel_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_23_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_368_obs_trg_cond , output \Core_2stage.DatPath_2stage.imm_z_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_0_obs_trg_cond , output core_io_interrupt_mtip_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._if_pc_next_T_7_obs_trg_cond , output \Core_2stage.DatPath_2stage._T_6_obs_trg_cond , output \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_19_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_15_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_tvm_obs_trg_cond , output \Core_2stage.c_io_ctl_mem_val_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_633_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_180_obs_trg_cond , output [2:0] \Core_2stage.DatPath_2stage._misaligned_mask_T_1_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_15_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_12_obs_trg_cond , output \Core_2stage.c_io_dmem_req_bits_fcn_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_46_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_3_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_13_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_ctl_if_kill_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_205_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_371_obs_trg_arg0 , output router_1_io_scratchPort_resp_valid_obs_trg_cond , output [10:0] \Core_2stage.DatPath_2stage._imm_j_sext_T_2_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mie_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_24_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_17_obs_trg_cond , output [4:0] \Core_2stage.DatPath_2stage.alu_shamt_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_8_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._bytes_T_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_1_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_31_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_192_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_25_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_1_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_scratchPort_resp_bits_data_obs_trg_cond , output [31:0] \SodorRequestRouter_2stage_1.io_corePort_req_bits_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_177_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_241_obs_trg_arg0 , output [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_mask_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_617_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_163_obs_trg_cond , output [2:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_req_bits_typ_obs_trg_arg0 , output \Core_2stage.d_io_ctl_exception_cause_obs_trg_cond , output [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_30_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_imem_req_bits_addr_state_invariant_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_dat_mem_store_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_183_obs_trg_arg0 , output \Core_2stage.d_io_dmem_req_bits_data_obs_trg_cond , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_107_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_3_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_288_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_0_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_95_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.if_pc_plus4_obs_trg_cond , output router_io_corePort_req_bits_data_obs_trg_cond , output [1:0] \Core_2stage.DatPath_2stage.csr_io_status_mpp_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_31_obs_trg_cond , output [2:0] \AsyncScratchPadMemory_2stage._io_core_ports_1_resp_bits_data_T_1_state_invariant_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_635_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_3_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_21_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_27_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_1_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_uxl_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_masterPort_req_bits_addr_obs_trg_cond , output io_master_port_1_resp_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_ube_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_3_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_addr_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_3_state_invariant_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_177_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_125_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.io_imem_resp_bits_data_state_invariant_obs_trg_arg0 , output [31:0] memory_io_debug_port_req_bits_addr_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_412_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._bytes_T_3_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_3_MPORT_en_obs_trg_cond , output \Core_2stage.DatPath_2stage.decode_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_19_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage._io_core_ports_1_resp_bits_data_T_1_state_invariant_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_192_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage.ctrl_pc_sel_obs_trg_arg0 , output [10:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._masks_mask_T_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_209_obs_trg_arg0 , output [2:0] io_debug_port_req_bits_typ_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_3_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_dmem_req_bits_typ_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_607_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_20_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_3_obs_trg_arg0 , output [7:0] \Core_2stage.DatPath_2stage._T_10_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_1_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.module_1_io_mem_data_0_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_622_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_15_obs_trg_cond , output \SodorRequestRouter_2stage_1.io_corePort_req_bits_addr_obs_trg_cond , output [31:0] router_io_masterPort_resp_bits_data_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_108_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_334_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_623_obs_trg_arg0 , output [11:0] \Core_2stage.DatPath_2stage.imm_s_obs_trg_arg0 , output [2:0] \SodorRequestRouter_2stage_0.io_corePort_req_bits_typ_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.cause_lsbs_obs_trg_cond , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1719_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mepc_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mpie_obs_trg_cond , output [32:0] \SodorRequestRouter_2stage_0._in_range_T_1_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_30_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_3_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.if_inst_buffer_valid_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_16_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_10_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_379_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_123_obs_trg_cond , output [31:0] \Core_2stage.d_io_imem_req_bits_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_csr_stall_obs_trg_arg0 , output \Core_2stage.d_io_dat_data_misaligned_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_0_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_1_obs_trg_cond , output \Core_2stage.c_io_ctl_exception_cause_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_wdata_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_corePort_req_valid_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_scratchPort_resp_valid_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_en_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_189_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_624_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_408_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_interrupt_T_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_11_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_corePort_resp_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_0_obs_trg_cond , output io_debug_port_req_valid_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_359_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._epc_T_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_242_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_363_obs_trg_arg0 , output [31:0] \Core_2stage.io_imem_resp_bits_data_state_invariant_obs_trg_arg0 , output [31:0] \Core_2stage.CtlPath_2stage.io_dat_inst_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.clock_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_631_obs_trg_cond , output \AsyncScratchPadMemory_2stage._io_core_ports_0_resp_bits_data_T_1_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_pc_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._GEN_1_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_272_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_3_MPORT_en_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_626_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_3_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_369_obs_trg_cond , output router_io_scratchPort_req_bits_fcn_obs_trg_arg0 , output [6:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_0_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_data_obs_trg_arg0 , output router_io_corePort_req_bits_fcn_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_289_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_325_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mtvec_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_12_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_595_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage.io_ctl_csr_cmd_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._bytes_T_3_obs_trg_cond , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_3_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_211_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_321_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.io_dmem_resp_bits_data_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_dat_csr_interrupt_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_1_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_365_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_20_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1714_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_77_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_wbdata_T_obs_trg_cond , output [62:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._shiftedVec_T_1_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_21_obs_trg_arg0 , output [7:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_zero1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.exe_reg_pc_obs_trg_cond , output \Core_2stage.DatPath_2stage._if_pc_next_T_3_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.if_pc_plus4_obs_trg_arg0 , output memory_io_core_ports_0_req_valid_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_125_obs_trg_arg0 , output [9:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_addr_state_invariant_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.module_1_io_mem_data_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_ctl_exception_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_dmem_resp_bits_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_0_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_594_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage._io_debug_port_resp_bits_data_T_1_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpv_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_corePort_req_bits_fcn_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_wbdata_T_2_obs_trg_cond , output \Core_2stage.io_interrupt_mtip_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._masks_maskWithOffset_T_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_time_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_26_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_arg0 , output [1:0] \Core_2stage.d_io_ctl_wb_sel_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_0_obs_trg_cond , output [20:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_addr_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_214_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.io_imem_resp_bits_data_state_invariant_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._imm_b_sext_T_2_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.exe_reg_inst_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_3_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_190_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_31_obs_trg_cond , output \Core_2stage.DatPath_2stage.imm_i_sext_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_interrupts_mtip_obs_trg_cond , output memory_io_core_ports_1_req_bits_addr_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_0_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_268_obs_trg_arg0 , output [62:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_19_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_18_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_tsr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_eret_obs_trg_arg0 , output \Core_2stage.c_io_ctl_rf_wen_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.csr_io_rw_wdata_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_size_obs_trg_arg0 , output \Core_2stage.d_reset_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.tval_inst_ma_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_13_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_upie_obs_trg_arg0 , output [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._large_r_T_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_zero1_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_mprv_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_266_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_316_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_jump_reg_target_T_1_obs_trg_cond , output router_io_respAddress_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_23_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_629_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_241_obs_trg_arg0 , output [6:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_op1_T_1_obs_trg_arg0 , output [31:0] \Core_2stage.io_imem_resp_bits_data_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_addr_obs_trg_cond , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.value_obs_trg_arg0 , output [9:0] \AsyncScratchPadMemory_2stage.mem_0_MPORT_addr_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_28_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_24_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_3_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_4_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_3_obs_trg_cond , output [31:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_data_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_18_obs_trg_arg0 , output \Core_2stage.d_io_ctl_if_kill_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.mem_0_MPORT_data_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_367_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_29_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_352_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_179_obs_trg_cond , output [5:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_34_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_124_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.addr_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_145_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.module__io_mem_data_0_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_mpie_obs_trg_cond , output io_debug_port_req_bits_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_108_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_8_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_368_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_rdata_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_620_obs_trg_cond , output [19:0] \Core_2stage.DatPath_2stage.imm_j_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._large_r_T_1_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_xs_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_cause_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_279_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.module_1_io_addr_obs_trg_cond , output \Core_2stage.c_io_imem_resp_valid_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.cs0_0_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mpie_obs_trg_arg0 , output [31:0] \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_data_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_0_MPORT_data_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_610_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_lo_lo_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.x86_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.offset_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_0_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._imm_i_sext_T_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_fs_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_539_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_182_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_0_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_12_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_283_obs_trg_arg0 , output [2:0] \Core_2stage.DatPath_2stage.io_ctl_csr_cmd_obs_trg_arg0 , output core_io_reset_vector_obs_trg_cond , output core_io_interrupt_meip_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_210_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_dat_mem_store_obs_trg_arg0 , output [1:0] \Core_2stage.d_io_ctl_op1_sel_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.module__io_mem_masks_3_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_12_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_3_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_3_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_122_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.debugTVec_obs_trg_cond , output [11:0] \Core_2stage.DatPath_2stage.csr_io_rw_addr_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_355_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_meip_obs_trg_cond , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1717_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_ungated_clock_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_89_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_3_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.module_1_io_mem_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_17_obs_trg_cond , output \SodorRequestRouter_2stage_0.io_respAddress_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_mtip_obs_trg_arg0 , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_3_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_269_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_600_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_2_MPORT_addr_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._io_dat_br_lt_T_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.exe_alu_out_obs_trg_cond , output [11:0] \Core_2stage.DatPath_2stage.imm_b_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_540_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_36_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugBreak_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_op1_T_4_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_67_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_exception_obs_trg_arg0 , output memory_io_core_ports_0_resp_valid_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_314_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.x79_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_310_obs_trg_cond , output \Core_2stage.DatPath_2stage._csr_io_tval_T_4_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_632_obs_trg_arg0 , output [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_13_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_5_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_isa_obs_trg_arg0 , output \Core_2stage.io_imem_req_bits_addr_state_invariant_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_wdata_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_115_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_msip_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_384_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugBreak_T_4_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_232_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_178_obs_trg_cond , output \SodorRequestRouter_2stage_0._in_range_T_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module_1_io_en_obs_trg_arg0 , output router_io_corePort_req_valid_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_0_obs_trg_cond , output \SodorRequestRouter_2stage_0.io_masterPort_resp_valid_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.sign_obs_trg_cond , output \Core_2stage.DatPath_2stage.imm_j_sext_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_26_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._csr_io_tval_T_6_obs_trg_arg0 , output [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_mask_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_MPORT_1_mask_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_31_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_1_MPORT_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_decode_0_read_illegal_T_16_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_5_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_ube_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_16_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_obs_trg_cond , output [19:0] \Core_2stage.DatPath_2stage._imm_s_sext_T_2_obs_trg_arg0 , output core_io_interrupt_debug_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_366_obs_trg_arg0 , output io_debug_port_req_bits_addr_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_ungated_clock_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_corePort_req_valid_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage.cs0_4_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_606_obs_trg_arg0 , output \Core_2stage.d_io_dat_data_misaligned_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_sd_rv32_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_339_obs_trg_arg0 , output memory_io_debug_port_req_bits_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_330_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_gva_obs_trg_cond , output \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_8_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_arg0 , output [9:0] \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.csr_io_pc_obs_trg_arg0 , output [4:0] \Core_2stage.DatPath_2stage.io_ctl_alu_fun_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_75_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_225_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_2_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._bytes_T_1_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_583_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_uie_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_364_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module__io_mem_masks_3_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_size_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._m_interrupts_T_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_mbe_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_debug_obs_trg_arg0 , output [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_maskWithOffset_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_221_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_217_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_11_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_618_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_4_obs_trg_cond , output \Core_2stage.d_io_dat_inst_misaligned_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tvm_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_175_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_2_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_246_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_128_obs_trg_cond , output [31:0] \AsyncScratchPadMemory_2stage.module__io_data_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage.io_ctl_mem_typ_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.exe_br_target_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_data_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.regfile_11_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_dat_if_valid_resp_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_1_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_interruptOffset_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_tval_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_25_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_239_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.anyInterrupt_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_29_obs_trg_cond , output \Core_2stage.DatPath_2stage.imm_i_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_322_obs_trg_cond , output \Core_2stage.d_io_reset_vector_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_10_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.wdata_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_ctl_op2_sel_obs_trg_cond , output [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_mask_obs_trg_arg0 , output \Core_2stage.c_io_dat_inst_obs_trg_cond , output [4:0] \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_addr_obs_trg_arg0 , output router_io_corePort_resp_valid_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_370_obs_trg_arg0 , output [15:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_7_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_uie_obs_trg_arg0 , output io_debug_port_req_bits_fcn_obs_trg_cond , output router_1_io_scratchPort_req_bits_typ_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.exe_br_target_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._bytes_T_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_0_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_dat_br_ltu_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.regfile_24_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_182_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_2_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_196_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_96_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.io_reset_vector_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_354_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._if_pc_next_T_2_obs_trg_cond , output router_1_io_scratchPort_req_valid_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_367_obs_trg_cond , output \SodorRequestRouter_2stage_0.io_corePort_req_valid_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_173_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_9_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_size_obs_trg_cond , output \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_fcn_obs_trg_arg0 , output [7:0] \Core_2stage.DatPath_2stage._T_8_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_7_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.sign_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_data_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_226_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.large__obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_102_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_op1_T_2_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_605_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_99_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_599_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage.io_ctl_wb_sel_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_op2_T_5_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_data_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_634_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_csr_stall_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_data_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_227_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sbe_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_masterPort_req_bits_typ_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_175_obs_trg_arg0 , output \Core_2stage.d_io_interrupt_meip_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_295_obs_trg_cond , output \SodorRequestRouter_2stage_0.io_corePort_resp_valid_obs_trg_cond , output router_io_masterPort_req_bits_fcn_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_332_obs_trg_cond , output \Core_2stage.DatPath_2stage._csr_io_tval_T_2_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_615_obs_trg_cond , output [2:0] core_io_dmem_req_bits_typ_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_117_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_49_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_98_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_165_obs_trg_arg0 , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_8_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_316_obs_trg_cond , output [31:0] router_io_scratchPort_req_bits_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_step_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_v_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._masks_maskWithOffset_T_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_28_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mstatus_T_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_interrupt_meip_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_signed_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_2_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_539_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_182_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_180_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_17_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_wbdata_T_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_mpp_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_interrupts_debug_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_interrupt_meip_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_3_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_628_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_293_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_11_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_mask_T_obs_trg_cond , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_218_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tsr_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._bytes_T_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_21_obs_trg_arg0 , output [9:0] \AsyncScratchPadMemory_2stage.mem_3_MPORT_addr_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_ctl_rf_wen_obs_trg_arg0 , output \Core_2stage.io_dmem_req_bits_typ_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_1_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_0_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_2_obs_trg_arg0 , output io_interrupt_debug_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_631_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_14_obs_trg_cond , output [6:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.nextSmall_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_53_obs_trg_arg0 , output [31:0] \Core_2stage.io_imem_req_bits_addr_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._masks_mask_T_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_8_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_393_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_dmem_req_bits_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_15_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_169_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_85_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_212_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_617_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_mask_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_390_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_data_obs_trg_arg0 , output \Core_2stage.c_io_ctl_pc_sel_obs_trg_cond , output \Core_2stage.DatPath_2stage._if_pc_next_T_1_obs_trg_arg0 , output [32:0] \SodorRequestRouter_2stage_1._resp_in_range_T_3_obs_trg_arg0 , output [9:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_addr_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.bytes_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._debugTVec_T_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_372_obs_trg_arg0 , output router_io_corePort_resp_bits_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_1_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_2_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_20_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_385_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_en_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.imm_j_sext_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.clock_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_signed_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_data_obs_trg_cond , output \Core_2stage.c_io_ctl_op2_sel_obs_trg_cond , output \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_debug_obs_trg_arg0 , output io_master_port_0_resp_bits_data_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_375_obs_trg_arg0 , output [31:0] io_master_port_1_req_bits_data_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_220_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_18_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_172_obs_trg_arg0 , output \Core_2stage.reset_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.system_insn_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._m_interrupts_T_5_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_12_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_3_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_212_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.exe_wbdata_obs_trg_arg0 , output [31:0] \SodorRequestRouter_2stage_0.io_corePort_req_bits_addr_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_cond , output [31:0] \Core_2stage.CtlPath_2stage.io_ctl_exception_cause_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_208_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_595_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_32_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_342_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_1_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_57_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_3_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_3_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_ungated_clock_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_15_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_16_obs_trg_cond , output \SodorRequestRouter_2stage_0.io_scratchPort_req_valid_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_31_obs_trg_arg0 , output \Core_2stage.d_io_ctl_stall_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_ctl_wb_sel_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.module_1_io_size_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mie_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.reg_interrupt_handled_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_367_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_35_obs_trg_arg0 , output [31:0] \SodorRequestRouter_2stage_0.io_scratchPort_resp_bits_data_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_65_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_376_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.wdata_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_285_obs_trg_cond , output [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_216_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_120_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_0_obs_trg_arg0 , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_19_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_19_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_1_obs_trg_cond , output \Core_2stage.c_io_dat_data_misaligned_obs_trg_cond , output \Core_2stage.d_io_dat_csr_eret_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_0_obs_trg_cond , output [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_71_obs_trg_cond , output io_master_port_0_req_valid_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_278_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_1_state_invariant_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_3_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_193_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_65_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._io_dat_data_misaligned_T_1_obs_trg_cond , output \Core_2stage.DatPath_2stage.reset_obs_trg_cond , output [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_2_obs_trg_arg0 , output \Core_2stage.io_imem_resp_valid_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_235_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_1_req_bits_addr_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_28_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_16_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_decode_0_read_illegal_T_16_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_334_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.clock_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_3_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_172_obs_trg_cond , output \Core_2stage.d_io_dat_csr_interrupt_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_105_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_173_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_117_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_op1_T_3_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.io_imem_req_bits_addr_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_2_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_19_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_313_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_corePort_req_bits_fcn_obs_trg_cond , output [31:0] io_master_port_1_resp_bits_data_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_dmem_req_valid_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_8_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_en_obs_trg_arg0 , output \Core_2stage.d_io_ctl_mem_val_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_393_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_uxl_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_215_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_1_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_ctl_csr_cmd_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_singleStep_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_383_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_mpie_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_11_obs_trg_cond , output \Core_2stage.d_io_dat_br_lt_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.io_imem_resp_bits_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._T_12_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_3_state_invariant_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_0_obs_trg_cond , output [20:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_addr_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_170_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_3_obs_trg_cond , output [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_hi_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_619_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_176_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_55_obs_trg_cond , output [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_214_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_26_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mie_obs_trg_arg0 , output \Core_2stage.d_io_dat_br_ltu_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_15_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.imm_j_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.io_dmem_req_bits_data_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_signed_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_MPORT_1_data_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_2_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_389_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_wbdata_T_6_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_217_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_fcn_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_1_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_374_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_331_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_corePort_req_bits_addr_obs_trg_cond , output \SodorRequestRouter_2stage_0.io_scratchPort_resp_bits_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_2_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_594_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_mask_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_79_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_3_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_108_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._shiftedVec_T_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_eret_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_1_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_271_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_op2_T_3_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_3_MPORT_addr_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_22_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_407_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_14_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_7_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.csr_io_status_isa_obs_trg_arg0 , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1714_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._sign_T_1_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_597_obs_trg_arg0 , output router_1_io_scratchPort_resp_bits_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_en_obs_trg_cond , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_12_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_1_obs_trg_arg0 , output router_io_masterPort_resp_valid_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_180_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_537_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_jump_reg_target_T_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_hi_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_ctl_mem_typ_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_op1_T_obs_trg_arg0 , output router_io_masterPort_req_bits_fcn_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_addr_obs_trg_cond , output [1:0] \Core_2stage.c_io_ctl_mem_fcn_obs_trg_arg0 , output io_interrupt_msip_obs_trg_cond , output [31:0] \Core_2stage.CtlPath_2stage._csignals_T_32_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_596_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_dmem_req_bits_fcn_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_603_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_79_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_1_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_283_obs_trg_cond , output [6:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_maskWithOffset_T_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_2_obs_trg_cond , output \Core_2stage.io_interrupt_debug_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_626_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_en_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_addr_state_invariant_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_176_obs_trg_cond , output [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_lo_obs_trg_arg0 , output [62:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._shiftedVec_T_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_108_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_3_obs_trg_cond , output \Core_2stage.io_interrupt_msip_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_289_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_12_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_0_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_18_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_typ_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_rw_cmd_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_540_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_13_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_25_obs_trg_arg0 , output memory_io_core_ports_1_resp_bits_data_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_dat_br_eq_obs_trg_cond , output \Core_2stage.DatPath_2stage._csr_io_tval_T_5_obs_trg_cond , output router_io_corePort_resp_valid_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_prv_obs_trg_arg0 , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_26_obs_trg_arg0 , output router_1_io_corePort_req_bits_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_59_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_sd_rv32_obs_trg_cond , output \Core_2stage.DatPath_2stage._T_1_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_310_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_214_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1722_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_5_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_addr_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_373_obs_trg_arg0 , output [31:0] \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_addr_obs_trg_arg0 , output \Core_2stage.d_io_dat_csr_eret_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_size_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_181_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_195_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_323_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_383_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_49_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_215_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_273_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_180_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpie_obs_trg_arg0 , output [32:0] \SodorRequestRouter_2stage_1._in_range_T_1_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_data_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_359_obs_trg_arg0 , output core_io_dmem_resp_valid_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_292_obs_trg_cond , output core_io_imem_resp_bits_data_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_622_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_15_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_290_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_corePort_resp_bits_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_doVector_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_3_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_dat_csr_eret_obs_trg_arg0 , output \Core_2stage.d_io_dat_csr_interrupt_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_7_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_signed_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_0_obs_trg_arg0 , output [10:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._masks_mask_T_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_3_obs_trg_cond , output router_1_io_corePort_req_valid_obs_trg_cond , output [31:0] router_io_respAddress_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_spie_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_616_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_380_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_data_obs_trg_arg0 , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_345_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_4_obs_trg_arg0 , output [31:0] router_1_io_masterPort_resp_bits_data_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_en_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_interrupt_msip_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_debug_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_dat_if_valid_resp_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_dat_csr_interrupt_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mip_obs_trg_cond , output \Core_2stage.c_io_ctl_mem_val_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_275_obs_trg_arg0 , output \Core_2stage.c_io_dat_if_valid_resp_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_wbdata_T_3_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_gva_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_195_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_18_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_2_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_ctl_exception_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._GEN_0_obs_trg_cond , output \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_15_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_637_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_214_obs_trg_cond , output [2:0] \Core_2stage.DatPath_2stage.io_ctl_op2_sel_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._bytes_T_1_obs_trg_cond , output [31:0] \SodorRequestRouter_2stage_1.io_masterPort_resp_bits_data_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_81_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_ctl_op1_sel_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_en_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_signed_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_1_obs_trg_arg0 , output [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_14_obs_trg_arg0 , output [31:0] \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_data_obs_trg_arg0 , output io_master_port_0_req_bits_typ_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_1_obs_trg_arg0 , output [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._masks_maskWithOffset_T_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_51_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_179_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_19_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_vs_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.sign_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_123_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_hi_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_336_obs_trg_cond , output [31:0] \AsyncScratchPadMemory_2stage.io_imem_req_bits_addr_state_invariant_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_102_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_corePort_resp_valid_obs_trg_arg0 , output [5:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_35_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_ctl_mem_fcn_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_23_obs_trg_arg0 , output router_io_scratchPort_req_bits_fcn_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_279_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_dat_inst_misaligned_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_2_state_invariant_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_312_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_287_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_274_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_21_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_1_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_184_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dpc_obs_trg_arg0 , output io_interrupt_debug_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_13_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage.io_dmem_req_bits_typ_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_masterPort_resp_valid_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_15_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_1_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_33_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_10_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_23_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_0_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_ctl_mem_fcn_obs_trg_cond , output core_io_imem_req_valid_obs_trg_cond , output memory_io_core_ports_0_req_bits_typ_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_28_obs_trg_arg0 , output router_io_scratchPort_resp_bits_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_37_obs_trg_cond , output \Core_2stage.c_io_dat_mem_store_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_sie_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_0_MPORT_mask_obs_trg_cond , output [31:0] router_io_corePort_resp_bits_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_296_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_12_obs_trg_cond , output \Core_2stage.DatPath_2stage._if_pc_next_T_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dpc_obs_trg_cond , output router_1_io_corePort_resp_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_MPORT_addr_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._sign_T_1_obs_trg_cond , output [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_73_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_interrupt_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_175_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_0_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_2_obs_trg_cond , output \Core_2stage.DatPath_2stage._if_pc_next_T_1_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._bytes_T_3_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_183_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.pending_interrupts_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_data_obs_trg_cond , output [1:0] \Core_2stage.DatPath_2stage.csr_io_status_prv_obs_trg_arg0 , output io_interrupt_meip_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_9_obs_trg_arg0 , output [31:0] \Core_2stage.io_imem_req_bits_addr_state_invariant_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_MPORT_data_obs_trg_arg0 , output [2:0] memory_io_core_ports_0_req_bits_typ_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_15_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_1_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_1_obs_trg_cond , output router_1_io_masterPort_req_bits_fcn_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_14_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_tvm_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.nextSmall_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_18_obs_trg_cond , output [6:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_interruptOffset_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_wbdata_T_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_dat_csr_interrupt_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_7_obs_trg_cond , output [20:0] \AsyncScratchPadMemory_2stage.module_1_io_addr_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_en_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_63_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_378_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_332_obs_trg_arg0 , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_14_obs_trg_arg0 , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_20_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.value_obs_trg_cond , output router_1_io_masterPort_req_valid_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_maskWithOffset_T_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_52_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_lo_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.exception_target_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_287_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_0_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_4_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_isa_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_ctl_rf_wen_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_99_obs_trg_cond , output core_io_imem_req_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.anyInterrupt_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_373_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_39_obs_trg_arg0 , output \Core_2stage.c_io_dmem_req_bits_fcn_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_masterPort_req_valid_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_19_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_fs_obs_trg_arg0 , output memory_io_core_ports_1_req_bits_typ_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_146_obs_trg_arg0 , output [31:0] \SodorRequestRouter_2stage_1.io_corePort_req_bits_data_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_285_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._bytes_T_3_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_data_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.regfile_18_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_281_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_224_obs_trg_cond , output memory_io_debug_port_req_bits_typ_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_168_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_0_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_6_obs_trg_cond , output \Core_2stage.d_io_ctl_stall_obs_trg_cond , output [82:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_hi_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_218_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_636_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugInt_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_20_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_2_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_3_obs_trg_arg0 , output \Core_2stage.io_imem_resp_valid_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_dat_data_misaligned_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mbe_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_0_MPORT_en_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_169_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_3_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_343_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_109_obs_trg_cond , output [4:0] \Core_2stage.CtlPath_2stage.rs1_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_cause_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_5_obs_trg_cond , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_115_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_1_obs_trg_cond , output [31:0] memory_io_core_ports_0_req_bits_data_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_masterPort_req_bits_fcn_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.pc_x_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_6_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_op1_T_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_48_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_41_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_signed_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_27_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_162_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_wfi_obs_trg_arg0 , output [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._large_r_T_3_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_obs_trg_cond , output [15:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mip_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_28_obs_trg_cond , output \SodorRequestRouter_2stage_0.io_corePort_req_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_24_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.if_reg_pc_obs_trg_arg0 , output io_imem_resp_bits_data_state_invariant_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_0_MPORT_addr_obs_trg_cond , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_318_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_1_MPORT_data_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_277_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_73_obs_trg_cond , output \Core_2stage.CtlPath_2stage.cs_val_inst_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_14_obs_trg_cond , output memory_io_core_ports_1_resp_valid_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_587_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_2_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_signed_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_2_MPORT_en_obs_trg_arg0 , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_34_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_interrupts_meip_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_mpv_obs_trg_cond , output [31:0] core_io_imem_req_bits_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_hartid_obs_trg_cond , output io_debug_port_resp_valid_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_197_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_174_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_609_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_call_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_en_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_320_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_cond , output \Core_2stage.CtlPath_2stage.cs0_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_11_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._sign_T_1_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_57_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_addr_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_380_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_24_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_data_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_387_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.tvec_obs_trg_cond , output [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_lo_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_retire_obs_trg_cond , output \Core_2stage.c_io_dat_inst_misaligned_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_debug_port_req_valid_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_103_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.exe_rs2_addr_obs_trg_cond , output [31:0] \Core_2stage.c_io_ctl_exception_cause_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._T_5_obs_trg_cond , output \Core_2stage.DatPath_2stage.imm_b_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_wfi_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_5_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.csr_wen_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_601_obs_trg_cond , output io_master_port_1_req_bits_data_obs_trg_cond , output [62:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._GEN_0_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_340_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_51_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_186_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_207_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_19_obs_trg_arg0 , output io_master_port_1_req_valid_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_311_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_meip_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_uie_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_MPORT_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_215_obs_trg_arg0 , output \Core_2stage.d_io_interrupt_debug_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_1_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_176_obs_trg_cond , output [5:0] \Core_2stage.DatPath_2stage._misaligned_mask_T_4_obs_trg_arg0 , output core_io_imem_resp_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_367_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_2_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_219_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage._T_14_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_293_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_spp_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_598_obs_trg_cond , output \Core_2stage.c_io_dat_csr_eret_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_3_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_26_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_344_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.exe_jump_reg_target_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_0_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._m_interrupts_T_3_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_2_obs_trg_cond , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.new_dcsr_ebreakm_obs_trg_arg0 , output [9:0] \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_arg0 , output core_clock_obs_trg_cond , output io_master_port_0_req_bits_fcn_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_634_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_48_obs_trg_cond , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_296_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_218_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_addr_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_1_req_valid_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_signed_obs_trg_arg0 , output io_debug_port_req_bits_fcn_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_187_obs_trg_arg0 , output [62:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._GEN_0_obs_trg_arg0 , output router_1_io_masterPort_req_bits_data_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.mem_2_MPORT_addr_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_47_obs_trg_cond , output [31:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_wfi_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_2_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_33_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_addr_obs_trg_arg0 , output \Core_2stage.d_io_dat_br_eq_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_206_obs_trg_arg0 , output [4:0] \Core_2stage.DatPath_2stage.exe_wbaddr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_op1_T_2_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_size_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_317_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_40_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupt_cause_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_wbdata_T_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_27_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.module_1_io_mem_addr_obs_trg_arg0 , output [31:0] \Core_2stage.CtlPath_2stage._csignals_T_38_obs_trg_arg0 , output \SodorRequestRouter_2stage_0._in_range_T_obs_trg_cond , output [31:0] router_1_io_scratchPort_req_bits_data_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_24_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_mxr_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.module_1_io_mem_data_3_obs_trg_cond , output [31:0] INSTR_inv_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_317_obs_trg_cond , output \Core_2stage.DatPath_2stage.clock_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_ebreakm_obs_trg_arg0 , output core_io_dmem_resp_bits_data_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_39_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_evec_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sie_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_1_obs_trg_cond , output core_reset_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_3_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_89_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_eret_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_244_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugTrigger_obs_trg_cond , output [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._masks_maskWithOffset_T_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.in_range_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_235_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_wbdata_T_5_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_1_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_316_obs_trg_cond , output \Core_2stage.d_io_imem_resp_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_95_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_0_MPORT_en_obs_trg_cond , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_100_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_33_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_ctl_mem_val_obs_trg_cond , output \Core_2stage.CtlPath_2stage.stall_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_115_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_dprv_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_231_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_dat_inst_misaligned_obs_trg_cond , output \SodorRequestRouter_2stage_0.io_masterPort_resp_bits_data_obs_trg_cond , output clock_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_338_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_22_obs_trg_cond , output \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_8_obs_trg_cond , output \Core_2stage.d_io_ctl_mem_fcn_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._bytes_T_1_obs_trg_arg0 , output [9:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_addr_obs_trg_arg0 , output [9:0] \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_addr_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_124_obs_trg_arg0 , output \Core_2stage.c_io_dat_br_ltu_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_377_obs_trg_cond , output [2:0] \SodorRequestRouter_2stage_1.io_masterPort_req_bits_typ_obs_trg_arg0 , output \Core_2stage.d_io_interrupt_msip_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_185_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_104_obs_trg_cond , output \Core_2stage.DatPath_2stage._if_pc_next_T_4_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_3_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_116_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_0_req_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_213_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_2_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_1_obs_trg_cond , output [31:0] \Core_2stage.c_io_dat_inst_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.misaligned_mask_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_7_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_29_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mcause_T_obs_trg_cond , output \SodorRequestRouter_2stage_0.io_scratchPort_req_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.exe_jmp_target_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_361_obs_trg_arg0 , output \Core_2stage.d_io_imem_req_valid_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_2_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dscratch_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_1_obs_trg_arg0 , output [4:0] \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_addr_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_15_obs_trg_cond , output [1:0] \Core_2stage.d_io_ctl_mem_fcn_obs_trg_arg0 , output \Core_2stage.io_dmem_req_valid_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_211_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_3_MPORT_mask_obs_trg_arg0 , output io_interrupt_meip_obs_trg_cond , output \Core_2stage.d_clock_obs_trg_cond , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_123_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_181_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_183_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_308_obs_trg_cond , output io_debug_port_req_bits_typ_obs_trg_cond , output [22:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_zero2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_cmd_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_318_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_lo_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_3_obs_trg_cond , output \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_12_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_319_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_3_obs_trg_cond , output [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_119_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_ctl_rf_wen_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_1_obs_trg_cond , output memory_io_core_ports_1_req_valid_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._bytes_T_3_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_ctl_pc_sel_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tvm_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_600_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_46_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_589_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_91_obs_trg_arg0 , output [19:0] \Core_2stage.DatPath_2stage.imm_u_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_3_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_239_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.clock_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_2_obs_trg_arg0 , output core_io_hartid_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._shiftedVec_T_1_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.module_1_io_mem_data_0_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_6_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_34_obs_trg_arg0 , output [2:0] \Core_2stage.DatPath_2stage.misaligned_mask_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_9_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_184_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_130_obs_trg_arg0 , output \Core_2stage.d_io_ctl_op2_sel_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_611_obs_trg_arg0 , output \Core_2stage.d_io_ctl_mem_val_obs_trg_arg0 , output core_io_dmem_req_valid_obs_trg_cond , output [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_xs_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_op2_T_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_83_obs_trg_arg0 , output [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_6_obs_trg_arg0 , output memory_clock_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_178_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_v_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_28_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_588_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_op2_T_4_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_246_obs_trg_cond , output [31:0] memory_io_debug_port_resp_bits_data_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_409_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_3_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_5_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_dprv_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_586_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_cease_obs_trg_cond , output [31:0] \SodorRequestRouter_2stage_0._resp_in_range_T_obs_trg_arg0 , output [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_cmd_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_6_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.io_dat_inst_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_1_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_326_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_7_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_45_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_debug_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_data_obs_trg_cond , output [20:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_addr_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_20_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_signed_obs_trg_cond , output \Core_2stage.DatPath_2stage.imm_u_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_93_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_imem_resp_bits_data_state_invariant_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_data_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_dat_mem_store_obs_trg_cond , output [2:0] router_io_corePort_req_bits_typ_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_389_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_407_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_2_MPORT_data_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_237_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_MPORT_1_en_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_3_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_0_state_invariant_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_182_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_35_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_sbe_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.imm_s_sext_obs_trg_arg0 , output router_1_io_respAddress_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease_r_obs_trg_cond , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_32_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_233_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._bytes_T_3_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_107_obs_trg_cond , output [7:0] \Core_2stage.DatPath_2stage.csr_io_status_zero1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_hartid_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_587_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_8_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_cond , output [2:0] \Core_2stage.c_io_ctl_pc_sel_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._sign_T_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_586_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_3_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_293_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._masks_mask_T_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reset_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_interrupt_msip_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_286_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_3_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_0_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_346_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_6_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_26_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_hie_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_3_obs_trg_cond , output memory_io_core_ports_0_resp_bits_data_obs_trg_cond , output [20:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_addr_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.module_1_io_data_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mie_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_621_obs_trg_arg0 , output memory_io_core_ports_0_req_bits_fcn_obs_trg_arg0 , output [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.large__obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_6_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_173_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_14_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sd_rv32_obs_trg_cond , output [1:0] \Core_2stage.DatPath_2stage.io_ctl_mem_fcn_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_118_obs_trg_arg0 , output [31:0] \SodorRequestRouter_2stage_1.io_scratchPort_resp_bits_data_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_101_obs_trg_arg0 , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_346_obs_trg_arg0 , output [31:0] memory_io_core_ports_1_req_bits_addr_obs_trg_arg0 , output \Core_2stage.d_io_ctl_alu_fun_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_343_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage.csr_cmd_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.imm_b_sext_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_ctl_if_kill_r_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_wfi_obs_trg_cond , output \Core_2stage.DatPath_2stage._GEN_11_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_356_obs_trg_cond , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_358_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._if_pc_next_T_4_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_0_obs_trg_cond , output \Core_2stage.DatPath_2stage._T_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_24_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_wfi_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_size_obs_trg_cond , output \Core_2stage.io_imem_req_bits_addr_obs_trg_cond , output [31:0] core_io_imem_resp_bits_data_obs_trg_arg0 , output [9:0] \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_327_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_303_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_305_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_spp_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_61_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugTrigger_T_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.imm_s_sext_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_ungated_clock_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_20_obs_trg_arg0 , output router_io_masterPort_req_valid_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_26_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_2_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_0_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_368_obs_trg_cond , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_111_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_op1_T_1_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.s_offset_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_335_obs_trg_arg0 , output [4:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._shiftedVec_T_obs_trg_arg0 , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_214_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_rw_addr_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.s_offset_obs_trg_cond , output [31:0] router_1_io_corePort_req_bits_data_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_186_obs_trg_cond , output \Core_2stage.CtlPath_2stage.cs0_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_342_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_294_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.csr_io_time_obs_trg_arg0 , output router_1_io_masterPort_req_bits_addr_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_fcn_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_10_obs_trg_cond , output core_io_dmem_req_bits_fcn_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_1_req_valid_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.s_offset_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_25_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_303_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_629_obs_trg_arg0 , output \Core_2stage.d_io_ctl_rf_wen_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_dat_br_eq_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_408_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_197_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_22_obs_trg_arg0 , output [5:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.small_1_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_18_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_ctl_if_kill_obs_trg_cond , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_36_obs_trg_arg0 , output \Core_2stage.c_io_dmem_resp_valid_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_300_obs_trg_cond , output [2:0] \Core_2stage.io_dmem_req_bits_typ_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.module_1_io_mem_data_2_obs_trg_cond , output \Core_2stage.c_io_dat_br_eq_obs_trg_cond , output \Core_2stage.DatPath_2stage._io_dat_br_lt_T_1_obs_trg_cond , output [31:0] \Core_2stage.d_io_dat_inst_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_97_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_uie_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_en_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.large_1_obs_trg_cond , output [31:0] RDATA_inv_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_2_obs_trg_cond , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_316_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_28_obs_trg_arg0 , output [62:0] \Core_2stage.DatPath_2stage._GEN_11_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_7_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_2_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_392_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_spp_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_193_obs_trg_cond , output [31:0] \SodorRequestRouter_2stage_0.io_respAddress_obs_trg_arg0 , output [6:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._GEN_1_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_data_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_cond , output [10:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._masks_mask_T_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.resp_in_range_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_117_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_dat_csr_eret_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._GEN_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_3_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_0_MPORT_mask_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_dprv_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.csr_io_status_vs_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_29_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_ctl_stall_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.offset_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_352_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_ctl_op1_sel_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_signed_state_invariant_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.value_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_1_obs_trg_cond , output \Core_2stage.DatPath_2stage._csr_io_tval_T_obs_trg_cond , output \Core_2stage.DatPath_2stage.imm_b_sext_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_240_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sbe_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_op2_T_4_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_35_obs_trg_cond , output [2:0] \AsyncScratchPadMemory_2stage._io_core_ports_0_resp_bits_data_T_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_99_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_hartid_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_2_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_609_obs_trg_cond , output router_io_scratchPort_req_valid_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_addr_obs_trg_cond , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.value_1_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_314_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_10_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_size_obs_trg_cond , output \Core_2stage.c_io_dat_if_valid_resp_obs_trg_cond , output io_master_port_1_req_bits_typ_obs_trg_cond , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_119_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_8_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_211_obs_trg_cond , output memory_io_core_ports_0_req_bits_fcn_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_size_obs_trg_cond , output \Core_2stage.c_io_dat_csr_interrupt_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_corePort_req_bits_typ_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_hartid_obs_trg_cond , output \SodorRequestRouter_2stage_0.io_masterPort_resp_valid_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_613_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_23_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_mbe_obs_trg_arg0 , output \Core_2stage.io_hartid_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_304_obs_trg_cond , output [31:0] memory_io_core_ports_1_resp_bits_data_obs_trg_arg0 , output \Core_2stage.c_io_dat_br_lt_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_dat_br_ltu_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_390_obs_trg_cond , output [2:0] \Core_2stage.DatPath_2stage.io_ctl_pc_sel_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcountinhibit_obs_trg_cond , output [31:0] \Core_2stage.io_dmem_req_bits_data_obs_trg_arg0 , output \Core_2stage.d_io_dat_if_valid_resp_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_masterPort_req_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_mie_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_607_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_maskWithOffset_obs_trg_cond , output router_1_io_masterPort_req_bits_typ_obs_trg_cond , output \Core_2stage.CtlPath_2stage.stall_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_hartid_obs_trg_cond , output router_io_corePort_req_bits_fcn_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.if_inst_buffer_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_116_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_410_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_en_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tw_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_215_obs_trg_arg0 , output [4:0] \Core_2stage.c_io_ctl_alu_fun_obs_trg_arg0 , output [104:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._new_mstatus_WIRE_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_274_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_602_obs_trg_arg0 , output [2:0] memory_io_debug_port_req_bits_typ_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_valid_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_122_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_27_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_269_obs_trg_arg0 , output memory_io_debug_port_resp_valid_obs_trg_cond , output [4:0] \Core_2stage.DatPath_2stage.exe_rs1_addr_obs_trg_arg0 , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_1_obs_trg_arg0 , output \Core_2stage.io_imem_resp_bits_data_state_invariant_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_232_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.sign_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_2_MPORT_en_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_194_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_data_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_343_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_14_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_633_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_3_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_dat_inst_misaligned_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_26_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_126_obs_trg_arg0 , output [31:0] io_master_port_0_req_bits_data_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_op2_T_6_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.exe_wbaddr_obs_trg_cond , output core_io_dmem_resp_valid_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage.io_ctl_op1_sel_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_18_obs_trg_cond , output io_master_port_0_resp_valid_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_ctl_rf_wen_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_25_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_96_obs_trg_arg0 , output \Core_2stage.c_io_imem_resp_valid_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_323_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_mask_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_wfi_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_309_obs_trg_arg0 , output [31:0] \Core_2stage.d_io_dmem_req_bits_addr_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_3_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_0_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_388_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_cond , output \Core_2stage.DatPath_2stage._tval_inst_ma_T_4_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_3_obs_trg_arg0 , output \Core_2stage.d_io_dat_inst_misaligned_obs_trg_arg0 , output [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_cause_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_hi_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease_r_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_230_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_597_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_imem_resp_bits_data_obs_trg_cond , output \Core_2stage.d_io_dat_br_ltu_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_28_obs_trg_cond , output [31:0] \SodorRequestRouter_2stage_1.io_corePort_resp_bits_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_8_obs_trg_cond , output [31:0] \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_addr_obs_trg_arg0 , output \Core_2stage.c_io_ctl_rf_wen_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_2_obs_trg_cond , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_122_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_276_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_imem_req_valid_obs_trg_arg0 , output \Core_2stage.d_io_interrupt_mtip_obs_trg_cond , output router_io_scratchPort_req_bits_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_op2_T_2_obs_trg_arg0 , output [31:0] \Core_2stage.d_io_ctl_exception_cause_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_data_obs_trg_cond , output [64:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_hi_hi_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_debug_port_resp_valid_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_7_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_upie_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_276_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_538_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_3_MPORT_data_obs_trg_cond , output \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_7_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._masks_maskWithOffset_T_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_sxl_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.offset_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_212_obs_trg_cond , output [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.large_1_obs_trg_arg0 , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_1_obs_trg_arg0 , output [2:0] \Core_2stage.DatPath_2stage.csr_io_rw_cmd_obs_trg_arg0 , output \SodorRequestRouter_2stage_0._resp_in_range_T_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_194_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_imem_resp_valid_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_18_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_reset_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_retire_obs_trg_arg0 , output core_io_interrupt_debug_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_1_obs_trg_cond , output \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_typ_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_16_obs_trg_cond , output \Core_2stage.c_io_dat_br_ltu_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.io_imem_req_bits_addr_state_invariant_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_19_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_174_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_0_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._io_dat_br_lt_T_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_73_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_10_obs_trg_cond , output io_master_port_1_req_valid_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_229_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_16_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_2_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_272_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_118_obs_trg_cond , output \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_11_obs_trg_cond , output \SodorRequestRouter_2stage_1._in_range_T_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_176_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_282_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_306_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_43_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugInt_T_1_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_97_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_11_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_32_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._bytes_T_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_spp_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_166_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_73_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_2_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_4_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._sign_T_1_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_207_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_36_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_vs_obs_trg_cond , output [2:0] \Core_2stage.c_io_dmem_req_bits_typ_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_2_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_cond , output [31:0] router_1_io_corePort_resp_bits_data_obs_trg_arg0 , output [1:0] \Core_2stage.c_io_ctl_op1_sel_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_69_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_374_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_0_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_120_obs_trg_cond , output memory_io_core_ports_0_req_bits_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_2_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module__io_addr_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module__io_mem_masks_2_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_3_obs_trg_arg0 , output [3:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_mask_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_282_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_176_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_ctl_exception_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_1_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.epc_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sum_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.bytes_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_MPORT_mask_obs_trg_cond , output \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_7_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_dmem_resp_valid_obs_trg_cond , output \Core_2stage.c_io_ctl_csr_cmd_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_188_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_15_obs_trg_arg0 , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_18_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_0_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_23_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_2_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_612_obs_trg_cond , output \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_fcn_obs_trg_cond , output \Core_2stage.c_io_ctl_exception_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_29_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_xs_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_270_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.bytes_obs_trg_cond , output \SodorRequestRouter_2stage_1._resp_in_range_T_1_obs_trg_cond , output [2:0] \Core_2stage.d_io_ctl_pc_sel_no_xept_obs_trg_arg0 , output [4:0] \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_addr_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_3_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_206_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_data_obs_trg_arg0 , output [7:0] \Core_2stage.DatPath_2stage._T_12_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_613_obs_trg_arg0 , output core_io_interrupt_meip_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_dat_data_misaligned_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.exception_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_19_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_183_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.m_interrupts_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_2_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_dat_br_ltu_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_437_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_sum_obs_trg_arg0 , output [20:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_addr_state_invariant_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_23_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcause_obs_trg_cond , output \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_22_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_12_obs_trg_cond , output \Core_2stage.c_io_ctl_exception_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_13_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_3_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_singleStepped_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_ctl_exception_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_18_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_23_obs_trg_arg0 , output \Core_2stage.io_dmem_req_bits_fcn_obs_trg_arg0 , output router_1_io_corePort_req_bits_fcn_obs_trg_arg0 , output [31:0] router_io_scratchPort_req_bits_data_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_606_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_interrupt_mtip_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.csr_io_cause_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_4_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_mask_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_3_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_signed_obs_trg_arg0 , output \Core_2stage.io_imem_req_valid_obs_trg_arg0 , output core_reset_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_185_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_279_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_csr_stall_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_2_state_invariant_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._GEN_0_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_op2_T_6_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_610_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_0_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_4_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_2_obs_trg_cond , output core_io_dmem_req_bits_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_21_obs_trg_cond , output \Core_2stage.c_io_ctl_stall_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_23_obs_trg_cond , output \Core_2stage.io_dmem_resp_bits_data_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_371_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.trapToDebug_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_411_obs_trg_arg0 , output \Core_2stage.c_io_ctl_mem_fcn_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_368_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_584_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_15_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_interrupts_msip_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.small_1_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_tval_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_addr_obs_trg_cond , output [31:0] router_1_io_respAddress_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_182_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_377_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_dat_br_lt_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_obs_trg_arg0 , output [7:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.cause_lsbs_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_dmem_req_bits_addr_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_625_obs_trg_arg0 , output io_imem_req_bits_addr_state_invariant_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_366_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_207_obs_trg_cond , output \Core_2stage.DatPath_2stage.exe_alu_op2_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_4_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_6_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_3_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_324_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._T_10_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_31_obs_trg_cond , output [4:0] \Core_2stage.d_io_ctl_alu_fun_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_2_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_630_obs_trg_cond , output \Core_2stage.c_io_ctl_pc_sel_no_xept_obs_trg_cond , output \Core_2stage.DatPath_2stage.if_inst_buffer_valid_obs_trg_cond , output [31:0] \Core_2stage.io_reset_vector_obs_trg_arg0 , output \Core_2stage.d_reset_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_maskWithOffset_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_37_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_26_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_436_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mie_T_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_365_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_0_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_130_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_28_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._sign_T_1_obs_trg_arg0 , output [6:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_2_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._masks_mask_T_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module__io_mem_data_1_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_238_obs_trg_cond , output [31:0] \Core_2stage.d_io_imem_resp_bits_data_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage.ctrl_pc_sel_no_xept_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mxr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_267_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_3_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_en_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._bytes_T_3_obs_trg_cond , output \Core_2stage.CtlPath_2stage.cs0_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sd_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_307_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_signed_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_ebreakm_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_388_obs_trg_arg0 , output [2:0] \SodorRequestRouter_2stage_0.io_masterPort_req_bits_typ_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_3_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_121_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mscratch_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_dv_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_5_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_632_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_12_obs_trg_arg0 , output io_master_port_0_req_bits_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_tw_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_MPORT_en_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_imem_resp_valid_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_maskWithOffset_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_MPORT_en_obs_trg_arg0 , output [31:0] \Core_2stage.io_dmem_resp_bits_data_obs_trg_arg0 , output \Core_2stage.c_io_ctl_op1_sel_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_245_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._new_mstatus_WIRE_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_216_obs_trg_cond , output \Core_2stage.c_io_ctl_stall_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_1_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_361_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_dmem_req_bits_fcn_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_15_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.csr_io_status_dprv_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_debug_port_resp_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_12_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_11_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_13_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_280_obs_trg_arg0 , output io_interrupt_mtip_obs_trg_cond , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_30_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_3_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_219_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_218_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_625_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_31_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_mie_obs_trg_arg0 , output io_master_port_1_req_bits_addr_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_0_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_eret_T_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sxl_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_15_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_0_state_invariant_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_corePort_resp_bits_data_obs_trg_cond , output \Core_2stage.DatPath_2stage._if_pc_next_T_5_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_0_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_ret_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_hi_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_en_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_180_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_mxr_obs_trg_cond , output \Core_2stage.io_imem_req_valid_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_7_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_masterPort_resp_valid_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_addr_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_ctl_stall_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_12_obs_trg_cond , output \Core_2stage.DatPath_2stage._misaligned_mask_T_1_obs_trg_cond , output [31:0] \Core_2stage.d_io_reset_vector_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_15_obs_trg_arg0 , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.addr_obs_trg_arg0 , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_2_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_26_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_wbdata_T_5_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_341_obs_trg_arg0 , output [31:0] memory_io_core_ports_0_req_bits_addr_obs_trg_arg0 , output core_io_imem_req_bits_addr_obs_trg_cond , output \Core_2stage.c_io_dat_br_eq_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.module__io_size_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_dv_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.csr_wen_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_588_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_op2_T_3_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_437_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_537_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_2_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_213_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_174_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpp_obs_trg_arg0 , output \Core_2stage.io_interrupt_mtip_obs_trg_cond , output \SodorRequestRouter_2stage_1._in_range_T_3_obs_trg_cond , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_mask_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_2_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_26_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_129_obs_trg_cond , output \Core_2stage.d_io_dat_mem_store_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module__io_mem_masks_2_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_18_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_eret_T_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_3_MPORT_mask_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_arg0 , output \Core_2stage.d_io_hartid_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpp_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_379_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_309_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_618_obs_trg_cond , output io_master_port_1_req_bits_fcn_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_maskWithOffset_obs_trg_cond , output \Core_2stage.DatPath_2stage.decode_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_7_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_en_obs_trg_cond , output [2:0] \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_typ_obs_trg_arg0 , output [4:0] \Core_2stage.DatPath_2stage.regfile_MPORT_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._T_1_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_18_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_2_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_222_obs_trg_arg0 , output [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_lo_obs_trg_arg0 , output [31:0] \SodorRequestRouter_2stage_1._in_range_T_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_0_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_29_obs_trg_cond , output router_1_io_scratchPort_req_bits_fcn_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.exe_wbdata_obs_trg_cond , output [20:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_13_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_dat_inst_misaligned_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_ret_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_19_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_31_obs_trg_arg0 , output \SodorRequestRouter_2stage_0._resp_in_range_T_1_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_singleStep_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_637_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_21_obs_trg_arg0 , output [31:0] router_1_io_masterPort_req_bits_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_MPORT_1_en_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_addr_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_291_obs_trg_cond , output \SodorRequestRouter_2stage_0.io_scratchPort_resp_valid_obs_trg_cond , output [1:0] \Core_2stage.DatPath_2stage.csr_io_status_sxl_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_10_obs_trg_arg0 , output \Core_2stage.d_clock_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_164_obs_trg_arg0 , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_219_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_27_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_244_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_20_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_4_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module__io_mem_addr_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module__io_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_3_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_0_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_ctl_exception_cause_obs_trg_cond , output core_io_dmem_req_valid_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_37_obs_trg_arg0 , output [2:0] \Core_2stage.d_io_ctl_op2_sel_obs_trg_arg0 , output [31:0] io_master_port_1_req_bits_addr_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_1_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_7_obs_trg_cond , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_130_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_interrupt_debug_obs_trg_cond , output [2:0] \Core_2stage.c_io_ctl_op2_sel_obs_trg_arg0 , output \Core_2stage.c_io_dat_mem_store_obs_trg_cond , output memory_io_debug_port_req_valid_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.exe_rs2_data_obs_trg_arg0 , output router_1_io_scratchPort_req_bits_fcn_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_3_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_imem_req_bits_addr_state_invariant_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._cause_T_5_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_addr_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_35_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.csr_io_status_xs_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_2_obs_trg_arg0 , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1722_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_ctl_mem_val_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_10_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_1_req_bits_typ_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_interrupt_mtip_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.small__obs_trg_cond , output \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_2_obs_trg_cond , output \Core_2stage.DatPath_2stage._csr_io_tval_T_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_127_obs_trg_cond , output [2:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_typ_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_327_obs_trg_cond , output \Core_2stage.DatPath_2stage._csr_io_tval_T_1_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_11_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_15_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.pending_interrupts_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_20_obs_trg_cond , output [2:0] \SodorRequestRouter_2stage_1.io_corePort_req_bits_typ_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_41_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_imem_resp_bits_data_state_invariant_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_26_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_357_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.x86_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_interrupts_mtip_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_2_obs_trg_arg0 , output \Core_2stage.d_io_dat_mem_store_obs_trg_arg0 , output \Core_2stage.io_dmem_resp_valid_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_clock_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_spp_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_sie_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_1_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_336_obs_trg_arg0 , output [10:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._masks_mask_T_obs_trg_arg0 , output [9:0] \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_604_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_reset_vector_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_603_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_cause_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_608_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_118_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_362_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_1_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.exe_rs1_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._if_pc_next_T_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_11_obs_trg_cond , output \Core_2stage.io_dmem_req_bits_addr_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_321_obs_trg_arg0 , output router_io_scratchPort_resp_valid_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_size_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._sign_T_1_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_357_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_25_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_2_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_277_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_imem_resp_valid_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.csr_io_interrupt_cause_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_scratchPort_req_valid_obs_trg_cond , output [31:0] core_io_reset_vector_obs_trg_arg0 , output \Core_2stage.reset_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_273_obs_trg_arg0 , output core_io_interrupt_mtip_obs_trg_cond , output \Core_2stage.DatPath_2stage.exception_target_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._csr_io_tval_T_5_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_fcn_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_12_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_19_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_23_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._cause_T_5_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_189_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.module__io_mem_data_3_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_186_obs_trg_cond , output memory_io_debug_port_resp_valid_obs_trg_arg0 , output [20:0] \AsyncScratchPadMemory_2stage.module__io_addr_obs_trg_arg0 , output [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_hi_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_386_obs_trg_arg0 , output \Core_2stage.d_io_dmem_resp_bits_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_214_obs_trg_cond , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mip_T_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_2_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_MPORT_1_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_331_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_14_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_205_obs_trg_arg0 , output memory_clock_obs_trg_cond , output router_1_io_masterPort_resp_valid_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_addr_obs_trg_cond , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_99_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_MPORT_mask_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_22_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_360_obs_trg_cond , output router_io_corePort_req_bits_addr_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_19_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_130_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_23_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_7_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_en_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugInt_T_1_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_9_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_4_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_0_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.s_offset_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_1_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_cease_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_410_obs_trg_cond , output router_io_masterPort_resp_bits_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_lo_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_636_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_0_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_109_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_2_MPORT_mask_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_lo_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_386_obs_trg_cond , output [31:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_data_obs_trg_arg0 , output memory_io_core_ports_0_req_bits_addr_obs_trg_cond , output \Core_2stage.io_dmem_resp_valid_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_412_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_fs_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_hie_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_241_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_size_state_invariant_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_165_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_19_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_1_obs_trg_cond , output \Core_2stage.c_io_dat_csr_interrupt_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mepc_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.reset_obs_trg_arg0 , output \Core_2stage.d_io_ctl_pc_sel_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_333_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.module_1_io_mem_data_3_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_isa_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_7_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_100_obs_trg_cond , output router_io_corePort_req_valid_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_3_obs_trg_cond , output router_1_io_masterPort_resp_valid_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_211_obs_trg_arg0 , output io_debug_port_resp_valid_obs_trg_arg0 , output [4:0] \Core_2stage.CtlPath_2stage.io_ctl_alu_fun_obs_trg_arg0 , output router_1_io_scratchPort_req_bits_data_obs_trg_cond , output router_1_io_corePort_req_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_12_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_239_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_12_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_31_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_mask_obs_trg_cond , output [31:0] \AsyncScratchPadMemory_2stage.module_1_io_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._csr_io_tval_T_1_obs_trg_cond , output io_master_port_1_resp_bits_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_ctl_alu_fun_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_ctl_stall_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_0_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_319_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_358_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._notDebugTVec_T_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_627_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.exe_jmp_target_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_170_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_size_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_en_obs_trg_arg0 , output \Core_2stage.clock_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_245_obs_trg_arg0 , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_maskWithOffset_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_31_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_zero2_obs_trg_cond , output \Core_2stage.CtlPath_2stage.cs0_0_obs_trg_arg0 , output [4:0] \Core_2stage.DatPath_2stage.exe_rs2_addr_obs_trg_arg0 , output \SodorRequestRouter_2stage_1._resp_in_range_T_obs_trg_cond , output [2:0] memory_io_core_ports_1_req_bits_typ_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.cs_alu_fun_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module__io_mem_masks_0_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_363_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_op2_T_2_obs_trg_cond , output [2:0] \Core_2stage.d_io_ctl_csr_cmd_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_data_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_328_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_329_obs_trg_cond , output router_1_io_masterPort_req_valid_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_183_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_typ_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_en_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module__io_mem_masks_1_obs_trg_cond , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_106_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_14_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_ctl_if_kill_r_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_wbdata_T_4_obs_trg_cond , output \Core_2stage.DatPath_2stage.if_reg_pc_obs_trg_cond , output \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_3_obs_trg_cond , output [12:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_28_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_25_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_87_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_298_obs_trg_cond , output [31:0] router_io_corePort_req_bits_data_obs_trg_arg0 , output router_io_scratchPort_req_bits_data_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_5_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.resp_in_range_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_1_obs_trg_arg0 , output [2:0] router_1_io_corePort_req_bits_typ_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_222_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_328_obs_trg_cond , output router_io_masterPort_req_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_108_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_20_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_242_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_163_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._if_pc_next_T_2_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_224_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.exe_reg_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_36_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_18_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_21_obs_trg_arg0 , output memory_io_debug_port_req_bits_fcn_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_170_obs_trg_cond , output \Core_2stage.d_io_ctl_pc_sel_no_xept_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_1_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_10_obs_trg_arg0 , output \Core_2stage.c_io_dat_inst_misaligned_obs_trg_cond , output core_io_interrupt_msip_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_20_obs_trg_cond , output [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._T_4_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._GEN_3_obs_trg_cond , output \Core_2stage.CtlPath_2stage.illegal_obs_trg_arg0 , output [2:0] \Core_2stage.c_io_ctl_pc_sel_no_xept_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_28_obs_trg_arg0 , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_ctl_op2_sel_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_354_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.s_offset_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_170_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_sd_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_223_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_eret_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_size_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_120_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_maskWithOffset_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_27_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_308_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_93_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sie_obs_trg_arg0 , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_3_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_call_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_tw_obs_trg_cond , output core_clock_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_7_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_dat_inst_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_13_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_3_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_2_obs_trg_cond , output [31:0] io_master_port_0_resp_bits_data_obs_trg_arg0 , output [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcountinhibit_obs_trg_arg0 , output [19:0] \Core_2stage.DatPath_2stage._imm_i_sext_T_2_obs_trg_arg0 , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_344_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_dat_mem_store_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.s_offset_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_zero2_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._bytes_T_1_obs_trg_arg0 , output [31:0] \Core_2stage.CtlPath_2stage._csignals_T_16_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_5_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.ctrl_pc_sel_obs_trg_cond , output [31:0] \SodorRequestRouter_2stage_0.io_corePort_req_bits_data_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_23_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_fcn_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_tsr_obs_trg_cond , output \SodorRequestRouter_2stage_1.io_corePort_req_bits_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_101_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module__io_mem_data_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_time_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_dat_if_valid_resp_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_dat_csr_eret_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mcountinhibit_T_1_obs_trg_cond , output [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_218_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_cause_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_debug_obs_trg_cond , output \SodorRequestRouter_2stage_0.io_corePort_req_bits_data_obs_trg_cond , output [20:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_addr_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_216_obs_trg_arg0 , output \Core_2stage.clock_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_req_bits_addr_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_11_obs_trg_arg0 , output \Core_2stage.d_io_ctl_exception_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_6_obs_trg_cond , output \Core_2stage.DatPath_2stage._csr_io_tval_T_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_168_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._tval_inst_ma_T_3_obs_trg_arg0 , output [31:0] \Core_2stage.CtlPath_2stage._csignals_T_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_wfi_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_21_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_167_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_599_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_en_obs_trg_cond , output router_1_io_scratchPort_req_valid_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_372_obs_trg_cond , output \SodorRequestRouter_2stage_1.io_masterPort_req_valid_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_mask_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_608_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_122_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_119_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._exe_wbdata_T_6_obs_trg_arg0 , output \Core_2stage.d_io_dat_br_eq_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_145_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_11_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_5_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_mpv_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.csr_io_status_uxl_obs_trg_arg0 , output router_io_scratchPort_resp_valid_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_mask_obs_trg_cond , output \Core_2stage.DatPath_2stage._misaligned_mask_T_4_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_15_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_18_obs_trg_arg0 , output \Core_2stage.io_imem_resp_bits_data_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._sign_T_1_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_masterPort_req_valid_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_3_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_209_obs_trg_cond , output \Core_2stage.DatPath_2stage._tval_inst_ma_T_3_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_381_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_ctl_pc_sel_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_3_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_3_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_2_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_172_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_28_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_71_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.exe_alu_op1_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.reg_interrupt_handled_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_signed_obs_trg_arg0 , output [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_17_obs_trg_arg0 , output [2:0] \Core_2stage.c_io_ctl_csr_cmd_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_12_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_409_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_ctl_alu_fun_obs_trg_cond , output \Core_2stage.d_io_ctl_csr_cmd_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_0_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_singleStep_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_data_obs_trg_cond , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_dmem_req_valid_obs_trg_arg0 , output router_1_io_corePort_req_bits_fcn_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_3_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_119_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_213_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_183_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_385_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_imem_req_bits_addr_obs_trg_cond , output [11:0] \Core_2stage.DatPath_2stage.imm_i_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_15_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_166_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.exe_rs1_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_10_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_debug_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.d_interrupts_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_MPORT_1_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtval_obs_trg_cond , output \Core_2stage.io_interrupt_meip_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mprv_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_2_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_270_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_311_obs_trg_arg0 , output [10:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_mask_T_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_time_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_182_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_mask_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.cs_val_inst_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_dv_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_353_obs_trg_cond , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_118_obs_trg_arg0 , output [31:0] router_io_masterPort_req_bits_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_step_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_en_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_23_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_v_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_280_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_23_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_108_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_ctl_if_kill_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_7_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_valid_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_295_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_1_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_17_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.io_ctl_exception_cause_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.io_ctl_op1_sel_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_185_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_mask_T_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_122_obs_trg_cond , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugBreak_T_3_obs_trg_arg0 , output \Core_2stage.c_io_ctl_if_kill_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_338_obs_trg_cond , output [15:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mip_T_obs_trg_arg0 , output \Core_2stage.c_io_dmem_resp_valid_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_27_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_27_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_26_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_13_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_17_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_3_obs_trg_arg0 , output [7:0] \Core_2stage.DatPath_2stage._T_16_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_2_obs_trg_cond , output [31:0] \SodorRequestRouter_2stage_0.io_corePort_resp_bits_data_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_291_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.module_1_io_mem_data_1_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_177_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_55_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_addr_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.sign_obs_trg_arg0 , output [4:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._shiftedVec_T_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.mem_1_MPORT_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_121_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module__io_mem_data_0_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_105_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.bytes_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_369_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_124_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_103_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_32_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_mask_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module__io_en_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_1_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_120_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_1_MPORT_mask_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_18_obs_trg_arg0 , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_1_obs_trg_arg0 , output \Core_2stage.d_io_ctl_if_kill_obs_trg_cond , output \Core_2stage.CtlPath_2stage.cs_br_type_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_313_obs_trg_cond , output \Core_2stage.DatPath_2stage._if_pc_next_T_6_obs_trg_cond , output \Core_2stage.io_reset_vector_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.module__io_mem_data_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.nextSmall_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_83_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_233_obs_trg_arg0 , output [31:0] \SodorRequestRouter_2stage_0.io_masterPort_req_bits_data_obs_trg_arg0 , output [31:0] io_imem_req_bits_addr_state_invariant_obs_trg_arg0 , output [11:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.debugTVec_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_rw_wdata_obs_trg_cond , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_300_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage.cs_br_type_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sxl_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_242_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_171_obs_trg_arg0 , output [31:0] \Core_2stage.d_io_dmem_req_bits_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_hie_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_5_obs_trg_cond , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._csr_io_tval_T_4_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_356_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpie_obs_trg_cond , output [31:0] core_io_dmem_req_bits_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._if_pc_next_T_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_gva_obs_trg_cond , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_104_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage.cs_alu_fun_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupt_obs_trg_arg0 , output \Core_2stage.c_io_dat_data_misaligned_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_342_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.tvec_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_lo_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_dat_br_lt_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcause_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_masterPort_req_bits_fcn_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_290_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_zero1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_2_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_620_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.csr_cmd_obs_trg_cond , output router_1_io_corePort_req_bits_typ_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.if_inst_buffer_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sd_rv32_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_322_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_344_obs_trg_arg0 , output io_debug_port_req_valid_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_0_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_cease_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_gva_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sum_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_27_obs_trg_cond , output [31:0] \SodorRequestRouter_2stage_1.io_masterPort_req_bits_data_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_dat_br_eq_obs_trg_arg0 , output memory_io_core_ports_0_req_valid_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_2_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_11_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_294_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_10_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_3_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_47_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_5_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugInt_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_hartid_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._if_pc_next_T_6_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_8_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_size_obs_trg_cond , output \Core_2stage.io_interrupt_debug_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_217_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_585_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_3_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_191_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_438_obs_trg_cond , output \Core_2stage.d_io_ctl_rf_wen_obs_trg_cond , output memory_io_debug_port_req_bits_data_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_19_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_284_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_2_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_0_req_valid_obs_trg_cond , output router_1_io_scratchPort_resp_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._GEN_3_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_589_obs_trg_cond , output [22:0] \Core_2stage.DatPath_2stage.csr_io_status_zero2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.exe_wben_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_0_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_77_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_26_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_fcn_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_typ_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_212_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.cause_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.csr_io_rw_rdata_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_585_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_5_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_61_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.csr_io_evec_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.exception_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_interrupts_meip_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_2_obs_trg_cond , output memory_io_core_ports_1_req_valid_obs_trg_arg0 , output \Core_2stage.d_io_dmem_req_bits_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_91_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_1_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_11_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_6_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_5_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_18_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_172_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_9_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_2_obs_trg_cond , output [6:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_maskWithOffset_T_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_12_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_382_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_318_obs_trg_cond , output [2:0] \Core_2stage.DatPath_2stage._io_dat_data_misaligned_T_1_obs_trg_arg0 , output \Core_2stage.c_io_ctl_wb_sel_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.x79_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_wbdata_T_3_obs_trg_cond , output [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_2_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_0_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.sign_obs_trg_arg0 , output [9:0] \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.exe_wben_obs_trg_arg0 , output memory_io_core_ports_1_resp_valid_obs_trg_cond , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_3_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._epc_T_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_v_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.exe_reg_pc_plus4_obs_trg_cond , output reset_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_10_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_611_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugBreak_T_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mie_T_obs_trg_cond , output \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_20_obs_trg_cond , output \Core_2stage.DatPath_2stage._T_4_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_sd_obs_trg_cond , output \SodorRequestRouter_2stage_0.io_corePort_req_bits_fcn_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_ctl_pc_sel_no_xept_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_596_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_179_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_3_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_1_obs_trg_arg0 , output [9:0] \AsyncScratchPadMemory_2stage.mem_1_MPORT_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_dv_obs_trg_cond , output \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_addr_obs_trg_cond , output [31:0] router_io_masterPort_req_bits_addr_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.clock_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_23_obs_trg_cond , output [32:0] \SodorRequestRouter_2stage_1._resp_in_range_T_1_obs_trg_arg0 , output \Core_2stage.d_io_imem_resp_valid_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_624_obs_trg_arg0 , output [32:0] \SodorRequestRouter_2stage_0._resp_in_range_T_3_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_5_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_1_obs_trg_cond , output [2:0] \AsyncScratchPadMemory_2stage._io_core_ports_1_resp_bits_data_T_1_obs_trg_arg0 , output [2:0] router_io_scratchPort_req_bits_typ_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_85_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._T_22_obs_trg_arg0 , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_298_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_281_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_interruptVec_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_mprv_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_out_T_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_spp_obs_trg_cond , output [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_hi_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_343_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_320_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._T_17_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_344_obs_trg_cond , output [2:0] router_io_masterPort_req_bits_typ_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sd_obs_trg_cond , output [2:0] io_master_port_0_req_bits_typ_obs_trg_arg0 , output \Core_2stage.io_dmem_req_valid_obs_trg_arg0 , output router_io_scratchPort_req_bits_typ_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_605_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_5_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_362_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_341_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_2_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_wbdata_T_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_294_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_34_obs_trg_cond , output [31:0] io_debug_port_req_bits_data_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_scratchPort_resp_valid_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_15_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_69_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mcause_T_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_interrupt_obs_trg_arg0 , output io_master_port_0_req_bits_addr_obs_trg_cond , output router_io_masterPort_req_bits_data_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_28_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.module__io_size_obs_trg_arg0 , output reset_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_dat_csr_eret_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_217_obs_trg_cond , output [32:0] \SodorRequestRouter_2stage_1._in_range_T_3_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_116_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_614_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.exe_reg_pc_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_masterPort_req_bits_fcn_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_366_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_275_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_284_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_623_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_dat_br_ltu_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.new_dcsr_ebreakm_obs_trg_cond , output \Core_2stage.io_dmem_req_bits_fcn_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_15_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_21_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_0_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage._exe_alu_op1_T_4_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_345_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_en_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_242_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_interrupt_cause_obs_trg_cond , output \Core_2stage.DatPath_2stage.exe_rs2_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module_1_io_size_obs_trg_cond , output [31:0] \SodorRequestRouter_2stage_1._resp_in_range_T_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_306_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_size_state_invariant_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_236_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_436_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_18_obs_trg_cond , output \Core_2stage.d_io_imem_resp_bits_data_obs_trg_cond , output router_io_masterPort_req_bits_addr_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.regfile_9_obs_trg_arg0 , output [5:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.small__obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_prv_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._m_interrupts_T_5_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_6_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_16_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_corePort_resp_valid_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_MPORT_1_mask_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_interrupt_debug_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_3_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_318_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._csr_io_tval_T_6_obs_trg_cond , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_112_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_4_obs_trg_arg0 , output \Core_2stage.d_io_ctl_wb_sel_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mprv_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_113_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_8_obs_trg_arg0 , output io_reset_vector_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_30_obs_trg_cond , output \Core_2stage.DatPath_2stage.exe_reg_valid_obs_trg_cond , output [2:0] \Core_2stage.d_io_ctl_pc_sel_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_corePort_req_bits_typ_obs_trg_cond , output [2:0] router_1_io_masterPort_req_bits_typ_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_26_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_221_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.imm_u_sext_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_612_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_304_obs_trg_arg0 , output [10:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_mask_T_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_186_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_315_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_45_obs_trg_arg0 , output io_hartid_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_411_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_315_obs_trg_cond , output \Core_2stage.DatPath_2stage._io_dat_br_lt_T_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.regfile_10_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_127_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_4_obs_trg_cond , output [1:0] \Core_2stage.DatPath_2stage.io_ctl_wb_sel_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_3_obs_trg_arg0 , output [31:0] router_1_io_scratchPort_req_bits_addr_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_97_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.exe_alu_op2_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_11_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_210_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_interrupts_debug_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_spie_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_627_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_en_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_123_obs_trg_cond , output \Core_2stage.c_io_dat_csr_eret_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_341_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.cs0_1_obs_trg_cond , output \SodorRequestRouter_2stage_0.resp_in_range_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_81_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_635_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_0_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_13_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_19_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_13_obs_trg_cond , output [31:0] \SodorRequestRouter_2stage_1.io_respAddress_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.mem_3_MPORT_data_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_4_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.cs0_4_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.regfile_1_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_584_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_ube_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_38_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_95_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_evec_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_dat_data_misaligned_obs_trg_arg0 , output router_io_masterPort_req_bits_typ_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_singleStep_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_prv_obs_trg_cond , output \Core_2stage.d_io_interrupt_debug_obs_trg_arg0 , output [9:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_addr_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_370_obs_trg_cond , output [2:0] \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_typ_obs_trg_arg0 , output \SodorRequestRouter_2stage_0._in_range_T_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugTrigger_T_1_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_67_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.io_masterPort_resp_bits_data_obs_trg_cond , output [21:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_lo_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_0_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_op1_T_3_obs_trg_cond , output router_io_masterPort_resp_valid_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_op2_T_obs_trg_arg0 , output \Core_2stage.d_io_dat_if_valid_resp_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_315_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_124_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_75_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.whichInterrupt_obs_trg_cond , output \AsyncScratchPadMemory_2stage.module_1_io_en_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_638_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_164_obs_trg_cond , output \Core_2stage.CtlPath_2stage.io_ctl_if_kill_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_signed_state_invariant_obs_trg_arg0 , output \Core_2stage.d_io_ctl_mem_typ_obs_trg_cond , output \Core_2stage.d_io_imem_req_valid_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_392_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_27_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_207_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugTrigger_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage._io_core_ports_1_resp_bits_data_T_1_obs_trg_cond , output io_interrupt_mtip_obs_trg_arg0 , output router_1_io_corePort_resp_bits_data_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_219_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_dat_if_valid_resp_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_en_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_0_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.csr_io_tval_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_2_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_4_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.offset_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_2_obs_trg_cond , output [14:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.d_interrupts_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpv_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mxr_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_0_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_op2_T_5_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_342_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_14_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_174_obs_trg_cond , output [6:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._GEN_1_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_293_obs_trg_arg0 , output [31:0] \Core_2stage.d_io_dmem_resp_bits_data_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_addr_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_593_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage.io_ctl_mem_fcn_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_ctl_mem_typ_obs_trg_cond , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_maskWithOffset_obs_trg_arg0 , output [11:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_addr_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dscratch_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_231_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_239_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_interruptVec_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_11_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.regfile_14_obs_trg_cond , output \SodorRequestRouter_2stage_0.io_masterPort_req_bits_fcn_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_retire_obs_trg_cond , output \Core_2stage.DatPath_2stage._misaligned_mask_T_3_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.system_insn_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_278_obs_trg_arg0 , output [7:0] \Core_2stage.DatPath_2stage._T_5_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_en_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_223_obs_trg_arg0 , output \Core_2stage.io_hartid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_7_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_628_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_175_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_18_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_imem_req_valid_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_3_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_addr_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_179_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_98_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_1_obs_trg_cond , output [31:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_data_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_267_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_178_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_35_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_375_obs_trg_cond , output io_master_port_0_resp_valid_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_1_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_188_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_190_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.s_offset_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_mask_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.in_range_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_353_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_imem_resp_valid_obs_trg_cond , output \Core_2stage.CtlPath_2stage.ctrl_pc_sel_no_xept_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.bytes_obs_trg_arg0 , output [32:0] \SodorRequestRouter_2stage_0._resp_in_range_T_1_obs_trg_arg0 , output io_debug_port_resp_bits_data_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_376_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_115_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_3_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._notDebugTVec_T_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_1_MPORT_mask_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.io_pc_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_391_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_3_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_121_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_21_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_10_obs_trg_arg0 , output [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_2_obs_trg_arg0 , output [31:0] io_imem_resp_bits_data_state_invariant_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_340_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_387_obs_trg_cond , output [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1._masks_maskWithOffset_T_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_status_sbe_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.imm_u_sext_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_signed_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_271_obs_trg_cond , output [6:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.nextSmall_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_17_obs_trg_arg0 , output \Core_2stage.io_interrupt_meip_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_9_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_279_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.module__io_mem_data_1_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_maskWithOffset_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.bytes_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_238_obs_trg_arg0 , output [1:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_op2_T_1_obs_trg_cond , output io_master_port_1_req_bits_fcn_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_355_obs_trg_arg0 , output io_interrupt_msip_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_604_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1719_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_171_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_0_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_addr_state_invariant_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_366_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_330_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_27_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._T_16_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_maskWithOffset_T_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_630_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_ctl_stall_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_162_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_0_obs_trg_arg0 , output \SodorRequestRouter_2stage_1.in_range_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_2_MPORT_mask_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_data_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.module__io_mem_masks_1_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_9_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_234_obs_trg_cond , output \Core_2stage.d_io_interrupt_meip_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._exe_alu_out_T_10_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_364_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_274_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_rdata_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_243_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_3_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_312_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_602_obs_trg_cond , output \Core_2stage.c_io_ctl_alu_fun_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_229_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_mask_obs_trg_arg0 , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugBreak_T_4_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_23_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_2_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_1_MPORT_en_obs_trg_cond , output [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._masks_maskWithOffset_T_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_324_obs_trg_cond , output \Core_2stage.d_io_dat_inst_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_53_obs_trg_cond , output core_io_dmem_req_bits_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_en_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.csr_ren_obs_trg_cond , output \Core_2stage.DatPath_2stage.alu_shamt_obs_trg_cond , output \Core_2stage.DatPath_2stage._T_obs_trg_arg0 , output [2:0] router_1_io_scratchPort_req_bits_typ_obs_trg_arg0 , output [31:0] io_reset_vector_obs_trg_arg0 , output [8:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_lo_lo_obs_trg_arg0 , output \Core_2stage.d_io_ctl_op1_sel_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_41_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_5_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.csr_io_rw_rdata_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_241_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_cond , output router_1_io_corePort_resp_valid_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_18_obs_trg_cond , output [31:0] \Core_2stage.io_dmem_req_bits_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.new_mstatus_mie_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_8_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_191_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._imm_j_sext_T_2_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.regfile_17_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_391_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_273_obs_trg_cond , output [31:0] \SodorRequestRouter_2stage_0._in_range_T_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_ctl_mem_val_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_1_MPORT_en_obs_trg_arg0 , output [20:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.imm_s_obs_trg_cond , output \Core_2stage.DatPath_2stage._csr_io_tval_T_3_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_616_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_218_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupt_obs_trg_cond , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_1_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtvec_obs_trg_arg0 , output [31:0] router_io_scratchPort_resp_bits_data_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.exe_rs1_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.sign_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_ctl_mem_val_obs_trg_arg0 , output memory_io_debug_port_req_valid_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_mask_obs_trg_arg0 , output [11:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._debugTVec_T_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_107_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_273_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_37_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_28_obs_trg_cond , output \Core_2stage.d_io_interrupt_mtip_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_2_obs_trg_arg0 , output \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_11_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_1_obs_trg_cond , output [31:0] \SodorRequestRouter_2stage_0.io_masterPort_resp_bits_data_obs_trg_arg0 , output core_io_interrupt_msip_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_size_obs_trg_arg0 , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_337_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_19_obs_trg_arg0 , output [31:0] \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_2_obs_trg_cond , output core_io_dmem_req_bits_typ_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_15_obs_trg_arg0 , output [4:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_1_obs_trg_arg0 , output \Core_2stage.c_io_dat_br_lt_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_222_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_ctl_pc_sel_no_xept_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_31_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_obs_trg_cond , output core_io_imem_resp_valid_obs_trg_cond , output [3:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_95_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_226_obs_trg_arg0 , output [2:0] \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_20_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_msip_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.imm_z_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_17_obs_trg_cond , output core_io_dmem_req_bits_fcn_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_data_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._T_177_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._epc_T_1_obs_trg_cond , output \SodorRequestRouter_2stage_1.io_masterPort_req_bits_typ_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mie_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_305_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_227_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupt_cause_obs_trg_cond , output io_master_port_0_req_valid_obs_trg_arg0 , output memory_io_core_ports_0_resp_valid_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reset_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_3_obs_trg_cond , output [7:0] \Core_2stage.DatPath_2stage._T_6_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage._tval_inst_ma_T_4_obs_trg_arg0 , output core_io_hartid_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_33_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_addr_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_196_obs_trg_cond , output \Core_2stage.DatPath_2stage.regfile_28_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_debug_port_req_valid_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2._bytes_T_1_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.sign_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._io_interrupt_T_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_addr_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_107_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_240_obs_trg_cond , output [1:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_size_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_174_obs_trg_cond , output \SodorRequestRouter_2stage_1.io_scratchPort_req_valid_obs_trg_arg0 , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_129_obs_trg_arg0 , output memory_io_debug_port_resp_bits_data_obs_trg_cond , output \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_1_state_invariant_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_mask_obs_trg_cond , output \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_mask_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_329_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_0_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_3_obs_trg_arg0 , output io_hartid_obs_trg_cond , output [63:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_294_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.imm_i_sext_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_3_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.regfile_2_obs_trg_arg0 , output [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_3_obs_trg_arg0 , output \SodorRequestRouter_2stage_0.io_scratchPort_resp_valid_obs_trg_arg0 , output [1:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_1_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.m_interrupts_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_3_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._shiftedVec_T_1_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_288_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mtvec_obs_trg_cond , output \Core_2stage.DatPath_2stage.io_dat_br_lt_obs_trg_cond , output \Core_2stage.CtlPath_2stage.illegal_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage._csignals_T_638_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_41_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_evec_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_addr_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_addr_obs_trg_cond , output router_1_io_corePort_req_bits_data_obs_trg_cond , output [31:0] io_debug_port_resp_bits_data_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.io_dat_br_lt_obs_trg_arg0 , output clock_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.regfile_25_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtvec_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_20_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_signed_obs_trg_cond , output [3:0] \Core_2stage.CtlPath_2stage._csignals_T_180_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_220_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_230_obs_trg_cond , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_360_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_111_obs_trg_cond , output [2:0] \Core_2stage.CtlPath_2stage.io_ctl_pc_sel_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage.trapToDebug_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_io_status_sum_obs_trg_cond , output [9:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_addr_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_0_obs_trg_arg0 , output [2:0] \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_typ_obs_trg_arg0 , output [15:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_hi_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_ctl_exception_cause_obs_trg_cond , output \Core_2stage.DatPath_2stage._exe_alu_out_T_31_obs_trg_cond , output \Core_2stage.CtlPath_2stage._csignals_T_63_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.pc_x_obs_trg_cond , output \SodorRequestRouter_2stage_1._in_range_T_1_obs_trg_cond , output [3:0] \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_mask_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_11_obs_trg_cond , output \Core_2stage.DatPath_2stage.csr_clock_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_40_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_339_obs_trg_cond , output \Core_2stage.d_io_hartid_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_27_obs_trg_arg0 , output \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_51_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._masks_mask_T_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage.new_mstatus_mie_obs_trg_arg0 , output [7:0] \Core_2stage.DatPath_2stage._T_14_obs_trg_arg0 , output \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_cond , output [2:0] \Core_2stage.DatPath_2stage.io_ctl_pc_sel_no_xept_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_621_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_0_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage.io_ctl_wb_sel_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_4_obs_trg_cond , output \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_size_obs_trg_cond , output \Core_2stage.DatPath_2stage.CSRFile_2stage._epc_T_obs_trg_cond , output \Core_2stage.DatPath_2stage._T_8_obs_trg_cond , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mcountinhibit_T_1_obs_trg_arg0 , output [7:0] \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_11_obs_trg_arg0 , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtval_obs_trg_arg0 , output \Core_2stage.CtlPath_2stage._csignals_T_87_obs_trg_arg0 , output [1:0] \Core_2stage.CtlPath_2stage._csignals_T_208_obs_trg_arg0 , output [1:0] \Core_2stage.c_io_ctl_wb_sel_obs_trg_arg0 );
	assign RDATA_inv_obs_trg_cond = ( \Core_2stage.DatPath_2stage._exe_wbdata_T_1 ) && ( ! ( \Core_2stage.DatPath_2stage._exe_wbdata_T ) ) ;
	assign RDATA_inv_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_data ;
	assign INSTR_inv_obs_trg_cond = ( ! \Core_2stage.DatPath_2stage.io_ctl_if_kill_r ) ;
	assign INSTR_inv_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_reg_inst ;
	assign \Core_2stage.DatPath_2stage.regfile_0_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_0_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_0 ;
	assign \Core_2stage.DatPath_2stage.regfile_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_1 ;
	assign \Core_2stage.DatPath_2stage.regfile_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_2 ;
	assign \Core_2stage.DatPath_2stage.regfile_3_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_3_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_3 ;
	assign \Core_2stage.DatPath_2stage.regfile_4_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_4_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_4 ;
	assign \Core_2stage.DatPath_2stage.regfile_5_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_5_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_5 ;
	assign \Core_2stage.DatPath_2stage.regfile_6_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_6_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_6 ;
	assign \Core_2stage.DatPath_2stage.regfile_7_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_7_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_7 ;
	assign \Core_2stage.DatPath_2stage.regfile_8_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_8_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_8 ;
	assign \Core_2stage.DatPath_2stage.regfile_9_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_9_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_9 ;
	assign \Core_2stage.DatPath_2stage.regfile_10_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_10_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_10 ;
	assign \Core_2stage.DatPath_2stage.regfile_11_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_11_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_11 ;
	assign \Core_2stage.DatPath_2stage.regfile_12_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_12_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_12 ;
	assign \Core_2stage.DatPath_2stage.regfile_13_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_13_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_13 ;
	assign \Core_2stage.DatPath_2stage.regfile_14_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_14_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_14 ;
	assign \Core_2stage.DatPath_2stage.regfile_15_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_15_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_15 ;
	assign \Core_2stage.DatPath_2stage.regfile_16_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_16_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_16 ;
	assign \Core_2stage.DatPath_2stage.regfile_17_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_17_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_17 ;
	assign \Core_2stage.DatPath_2stage.regfile_18_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_18_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_18 ;
	assign \Core_2stage.DatPath_2stage.regfile_19_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_19_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_19 ;
	assign \Core_2stage.DatPath_2stage.regfile_20_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_20_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_20 ;
	assign \Core_2stage.DatPath_2stage.regfile_21_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_21_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_21 ;
	assign \Core_2stage.DatPath_2stage.regfile_22_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_22_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_22 ;
	assign \Core_2stage.DatPath_2stage.regfile_23_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_23_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_23 ;
	assign \Core_2stage.DatPath_2stage.regfile_24_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_24_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_24 ;
	assign \Core_2stage.DatPath_2stage.regfile_25_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_25_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_25 ;
	assign \Core_2stage.DatPath_2stage.regfile_26_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_26_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_26 ;
	assign \Core_2stage.DatPath_2stage.regfile_27_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_27_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_27 ;
	assign \Core_2stage.DatPath_2stage.regfile_28_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_28_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_28 ;
	assign \Core_2stage.DatPath_2stage.regfile_29_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_29_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_29 ;
	assign \Core_2stage.DatPath_2stage.regfile_30_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_30_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_30 ;
	assign \Core_2stage.DatPath_2stage.regfile_31_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_31_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_31 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._GEN_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._bytes_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._bytes_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._bytes_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._bytes_T_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._bytes_T_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._bytes_T_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_10_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_10_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_10 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_11_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_11_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_11 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_12_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_12_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_12 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_15_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_15_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_15 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_18_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_18_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_18 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_19_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_19_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_19 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_20_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_20_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_20 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_23_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_23_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_23 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_26_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_26_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_26 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_27_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_27_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_27 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_28_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_28_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_28 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_31_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_31_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_31 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_4_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_4_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_4 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_7_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_7_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._maskedVec_T_7 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._masks_maskWithOffset_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._masks_maskWithOffset_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._masks_maskWithOffset_T ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._masks_mask_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._masks_mask_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._masks_mask_T ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._shiftedVec_T_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._sign_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0._sign_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0._sign_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.bytes_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.bytes_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.bytes ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_addr ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_hi_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_hi_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_hi ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_lo_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_lo_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_data_lo ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_addr ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_mem_data_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_signed_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_signed_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_signed ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_size_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_size_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.io_size ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.maskedVec_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_mask_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_mask_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_mask ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_maskWithOffset_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_maskWithOffset_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.masks_maskWithOffset ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.s_offset_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.s_offset_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.s_offset ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.shiftedVec_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.sign_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_0.sign_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_0.sign ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._GEN_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._bytes_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._bytes_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._bytes_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._bytes_T_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._bytes_T_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._bytes_T_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_10_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_10_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_10 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_11_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_11_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_11 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_12_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_12_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_12 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_15_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_15_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_15 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_18_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_18_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_18 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_19_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_19_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_19 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_20_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_20_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_20 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_23_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_23_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_23 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_26_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_26_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_26 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_27_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_27_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_27 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_28_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_28_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_28 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_31_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_31_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_31 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_4_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_4_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_4 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_7_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_7_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._maskedVec_T_7 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._masks_maskWithOffset_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._masks_maskWithOffset_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._masks_maskWithOffset_T ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._masks_mask_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._masks_mask_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._masks_mask_T ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._shiftedVec_T_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._sign_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1._sign_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1._sign_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.bytes_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.bytes_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.bytes ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_addr ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_hi_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_hi_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_hi ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_lo_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_lo_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_data_lo ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_addr ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_mem_data_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_signed_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_signed_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_signed ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_size_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_size_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.io_size ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.maskedVec_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_mask_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_mask_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_mask ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_maskWithOffset_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_maskWithOffset_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.masks_maskWithOffset ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.s_offset_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.s_offset_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.s_offset ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.shiftedVec_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.sign_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_1.sign_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_1.sign ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._GEN_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._bytes_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._bytes_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._bytes_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._bytes_T_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._bytes_T_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._bytes_T_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_10_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_10_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_10 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_11_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_11_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_11 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_12_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_12_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_12 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_15_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_15_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_15 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_18_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_18_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_18 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_19_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_19_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_19 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_20_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_20_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_20 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_23_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_23_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_23 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_26_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_26_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_26 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_27_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_27_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_27 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_28_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_28_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_28 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_31_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_31_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_31 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_4_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_4_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_4 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_7_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_7_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._maskedVec_T_7 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._masks_maskWithOffset_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._masks_maskWithOffset_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._masks_maskWithOffset_T ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._masks_mask_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._masks_mask_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._masks_mask_T ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._shiftedVec_T_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._sign_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2._sign_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2._sign_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.bytes_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.bytes_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.bytes ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_addr ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_hi_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_hi_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_hi ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_lo_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_lo_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_data_lo ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_addr ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_mem_data_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_signed_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_signed_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_signed ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_size_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_size_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.io_size ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.maskedVec_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_mask_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_mask_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_mask ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_maskWithOffset_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_maskWithOffset_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.masks_maskWithOffset ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.s_offset_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.s_offset_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.s_offset ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.shiftedVec_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.sign_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_2.sign_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_2.sign ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._GEN_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._bytes_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._bytes_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._bytes_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._bytes_T_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._bytes_T_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._bytes_T_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_10_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_10_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_10 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_11_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_11_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_11 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_12_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_12_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_12 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_15_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_15_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_15 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_18_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_18_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_18 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_19_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_19_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_19 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_20_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_20_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_20 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_23_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_23_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_23 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_26_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_26_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_26 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_27_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_27_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_27 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_28_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_28_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_28 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_31_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_31_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_31 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_4_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_4_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_4 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_7_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_7_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._maskedVec_T_7 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._masks_maskWithOffset_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._masks_maskWithOffset_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._masks_maskWithOffset_T ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._masks_mask_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._masks_mask_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._masks_mask_T ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._shiftedVec_T_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._sign_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._sign_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant._sign_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.bytes_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.bytes_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.bytes ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_addr ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_hi_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_hi_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_hi ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_lo_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_lo_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_data_lo ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_addr ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_mem_data_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_signed_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_signed_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_signed ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_size_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_size_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.io_size ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.maskedVec_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_mask_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_mask_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_mask ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_maskWithOffset_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_maskWithOffset_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.masks_maskWithOffset ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.s_offset_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.s_offset_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.s_offset ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_0 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_2 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.shiftedVec_3 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.sign_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.sign_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemReader_2stage_state_invariant.sign ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._GEN_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._GEN_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._GEN_0 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._GEN_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._GEN_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._GEN_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_3 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_5_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_5_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_T_5 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_maskWithOffset_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_maskWithOffset_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_maskWithOffset_T ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_mask_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_mask_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._masks_mask_T ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._shiftedVec_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._shiftedVec_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._shiftedVec_T ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._shiftedVec_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._shiftedVec_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0._shiftedVec_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_addr ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_data ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_en ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_addr ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_0 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_2 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_data_3 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_0 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_2 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_mem_masks_3 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_size_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_size_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.io_size ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_0 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_2 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_3 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_mask_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_mask_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_mask ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_maskWithOffset_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_maskWithOffset_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.masks_maskWithOffset ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.offset_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.offset_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.offset ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_2 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_hi_3 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_2 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_0.shiftedVec_lo_3 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._GEN_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._GEN_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._GEN_0 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._GEN_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._GEN_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._GEN_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_3 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_5_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_5_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_T_5 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_maskWithOffset_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_maskWithOffset_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_maskWithOffset_T ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_mask_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_mask_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._masks_mask_T ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._shiftedVec_T_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._shiftedVec_T_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._shiftedVec_T ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._shiftedVec_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._shiftedVec_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1._shiftedVec_T_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_addr ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_data ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_en ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_addr ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_0 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_2 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_data_3 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_0 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_2 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_mem_masks_3 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_size_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_size_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.io_size ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_0 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_2 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_3 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_mask_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_mask_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_mask ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_maskWithOffset_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_maskWithOffset_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.masks_maskWithOffset ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.offset_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.offset_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.offset ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_2 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_hi_3 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_2 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.MemWriter_2stage_1.shiftedVec_lo_3 ;
	assign \AsyncScratchPadMemory_2stage._io_core_ports_0_resp_bits_data_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage._io_core_ports_0_resp_bits_data_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage._io_core_ports_0_resp_bits_data_T_1 ;
	assign \AsyncScratchPadMemory_2stage._io_core_ports_1_resp_bits_data_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage._io_core_ports_1_resp_bits_data_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage._io_core_ports_1_resp_bits_data_T_1 ;
	assign \AsyncScratchPadMemory_2stage._io_core_ports_1_resp_bits_data_T_1_state_invariant_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage._io_core_ports_1_resp_bits_data_T_1_state_invariant_obs_trg_arg0 = \AsyncScratchPadMemory_2stage._io_core_ports_1_resp_bits_data_T_1_state_invariant ;
	assign \AsyncScratchPadMemory_2stage._io_debug_port_resp_bits_data_T_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage._io_debug_port_resp_bits_data_T_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage._io_debug_port_resp_bits_data_T_1 ;
	assign \AsyncScratchPadMemory_2stage.clock_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.clock_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.clock ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_addr ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_data ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_fcn_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_fcn_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_fcn ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_typ_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_typ_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_req_bits_typ ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_req_valid_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_req_valid_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_req_valid ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_addr ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_data ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_addr ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_0 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_2 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_mem_data_3 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_signed_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_signed_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_signed ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_size_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_size_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_bits_data_module_io_size ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_valid_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_valid_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_0_resp_valid ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_req_bits_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_req_bits_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_req_bits_addr ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_req_bits_typ_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_req_bits_typ_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_req_bits_typ ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_req_valid_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_req_valid_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_req_valid ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_addr ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_addr_state_invariant_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_addr_state_invariant_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_addr_state_invariant ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_data ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_addr ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_addr_state_invariant_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_addr_state_invariant_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_addr_state_invariant ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_0 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_0_state_invariant_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_0_state_invariant_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_0_state_invariant ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_1_state_invariant_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_1_state_invariant_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_1_state_invariant ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_2 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_2_state_invariant_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_2_state_invariant_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_2_state_invariant ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_3 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_3_state_invariant_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_3_state_invariant_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_mem_data_3_state_invariant ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_signed_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_signed_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_signed ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_signed_state_invariant_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_signed_state_invariant_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_signed_state_invariant ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_size_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_size_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_size ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_size_state_invariant_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_size_state_invariant_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_bits_data_module_io_size_state_invariant ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_valid_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_valid_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_core_ports_1_resp_valid ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_addr ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_data ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_fcn_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_fcn_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_fcn ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_typ_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_typ_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_req_bits_typ ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_req_valid_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_req_valid_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_req_valid ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_addr ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_data ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_addr ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_0 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_2 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_mem_data_3 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_signed_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_signed_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_signed ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_size_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_size_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_resp_bits_data_module_io_size ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_valid_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_debug_port_resp_valid_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_debug_port_resp_valid ;
	assign \AsyncScratchPadMemory_2stage.io_imem_req_bits_addr_state_invariant_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_imem_req_bits_addr_state_invariant_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_imem_req_bits_addr_state_invariant ;
	assign \AsyncScratchPadMemory_2stage.io_imem_resp_bits_data_state_invariant_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.io_imem_resp_bits_data_state_invariant_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.io_imem_resp_bits_data_state_invariant ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_data ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_en ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_mask_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_mask_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_MPORT_1_mask ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_mask_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_MPORT_mask_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_MPORT_mask ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_0_resp_bits_data_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_io_core_ports_1_resp_bits_data_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_0_io_debug_port_resp_bits_data_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_data ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_en ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_mask_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_mask_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_MPORT_1_mask ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_mask_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_MPORT_mask_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_MPORT_mask ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_0_resp_bits_data_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_io_core_ports_1_resp_bits_data_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_1_io_debug_port_resp_bits_data_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_data ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_en ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_mask_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_mask_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_MPORT_1_mask ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_mask_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_MPORT_mask_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_MPORT_mask ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_0_resp_bits_data_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_io_core_ports_1_resp_bits_data_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_2_io_debug_port_resp_bits_data_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_data ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_en ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_mask_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_mask_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_MPORT_1_mask ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_mask_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_MPORT_mask_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_MPORT_mask ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_0_resp_bits_data_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_io_core_ports_1_resp_bits_data_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_addr ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_data ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.mem_3_io_debug_port_resp_bits_data_MPORT_en ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module_1_io_addr ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module_1_io_data ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module_1_io_en ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module_1_io_mem_addr ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_data_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_data_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module_1_io_mem_data_0 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_data_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_data_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module_1_io_mem_data_1 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_data_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_data_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module_1_io_mem_data_2 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_data_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_data_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module_1_io_mem_data_3 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_0 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_1 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_2 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module_1_io_mem_masks_3 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_size_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module_1_io_size_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module_1_io_size ;
	assign \AsyncScratchPadMemory_2stage.module__io_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module__io_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module__io_addr ;
	assign \AsyncScratchPadMemory_2stage.module__io_data_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module__io_data_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module__io_data ;
	assign \AsyncScratchPadMemory_2stage.module__io_en_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module__io_en_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module__io_en ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_addr_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_addr_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module__io_mem_addr ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_data_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_data_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module__io_mem_data_0 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_data_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_data_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module__io_mem_data_1 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_data_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_data_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module__io_mem_data_2 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_data_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_data_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module__io_mem_data_3 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_masks_0_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_masks_0_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module__io_mem_masks_0 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_masks_1_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_masks_1_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module__io_mem_masks_1 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_masks_2_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_masks_2_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module__io_mem_masks_2 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_masks_3_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module__io_mem_masks_3_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module__io_mem_masks_3 ;
	assign \AsyncScratchPadMemory_2stage.module__io_size_obs_trg_cond = 1 ;
	assign \AsyncScratchPadMemory_2stage.module__io_size_obs_trg_arg0 = \AsyncScratchPadMemory_2stage.module__io_size ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_1_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_11_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_11_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_11 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_13_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_13_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_13 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_130_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_130_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_130 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_15_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_15_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_15 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_16_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_16_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_16 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_162_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_162_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_162 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_163_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_163_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_163 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_164_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_164_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_164 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_165_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_165_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_165 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_166_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_166_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_166 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_167_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_167_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_167 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_168_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_168_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_168 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_169_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_169_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_169 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_17_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_17_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_17 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_170_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_170_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_170 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_171_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_171_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_171 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_172_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_172_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_172 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_173_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_173_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_173 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_174_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_174_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_174 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_175_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_175_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_175 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_176_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_176_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_176 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_177_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_177_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_177 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_178_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_178_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_178 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_179_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_179_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_179 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_180_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_180_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_180 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_181_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_181_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_181 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_182_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_182_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_182 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_183_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_183_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_183 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_184_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_184_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_184 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_185_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_185_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_185 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_186_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_186_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_186 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_187_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_187_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_187 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_188_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_188_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_188 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_189_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_189_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_189 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_19_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_19_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_19 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_190_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_190_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_190 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_191_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_191_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_191 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_192_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_192_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_192 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_193_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_193_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_193 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_194_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_194_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_194 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_195_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_195_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_195 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_196_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_196_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_196 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_197_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_197_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_197 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_205_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_205_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_205 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_206_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_206_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_206 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_207_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_207_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_207 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_208_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_208_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_208 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_209_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_209_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_209 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_21_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_21_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_21 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_210_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_210_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_210 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_211_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_211_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_211 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_212_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_212_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_212 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_213_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_213_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_213 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_214_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_214_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_214 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_215_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_215_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_215 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_216_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_216_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_216 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_217_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_217_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_217 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_218_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_218_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_218 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_219_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_219_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_219 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_220_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_220_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_220 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_221_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_221_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_221 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_222_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_222_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_222 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_223_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_223_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_223 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_224_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_224_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_224 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_225_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_225_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_225 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_226_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_226_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_226 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_227_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_227_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_227 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_228_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_228_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_228 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_229_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_229_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_229 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_23_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_23_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_23 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_230_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_230_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_230 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_231_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_231_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_231 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_232_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_232_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_232 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_233_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_233_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_233 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_234_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_234_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_234 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_235_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_235_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_235 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_236_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_236_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_236 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_237_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_237_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_237 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_238_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_238_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_238 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_239_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_239_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_239 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_240_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_240_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_240 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_241_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_241_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_241 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_242_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_242_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_242 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_243_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_243_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_243 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_244_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_244_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_244 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_245_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_245_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_245 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_246_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_246_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_246 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_25_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_25_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_25 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_266_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_266_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_266 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_267_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_267_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_267 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_268_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_268_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_268 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_269_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_269_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_269 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_27_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_27_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_27 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_270_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_270_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_270 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_271_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_271_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_271 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_272_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_272_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_272 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_273_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_273_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_273 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_274_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_274_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_274 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_275_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_275_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_275 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_276_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_276_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_276 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_277_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_277_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_277 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_278_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_278_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_278 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_279_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_279_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_279 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_280_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_280_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_280 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_281_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_281_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_281 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_282_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_282_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_282 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_283_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_283_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_283 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_284_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_284_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_284 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_285_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_285_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_285 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_286_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_286_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_286 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_287_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_287_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_287 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_288_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_288_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_288 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_289_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_289_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_289 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_29_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_29_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_29 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_290_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_290_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_290 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_291_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_291_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_291 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_292_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_292_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_292 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_293_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_293_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_293 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_294_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_294_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_294 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_295_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_295_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_295 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_3_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_3_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_3 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_303_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_303_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_303 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_304_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_304_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_304 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_305_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_305_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_305 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_306_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_306_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_306 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_307_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_307_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_307 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_308_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_308_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_308 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_309_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_309_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_309 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_31_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_31_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_31 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_310_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_310_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_310 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_311_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_311_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_311 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_312_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_312_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_312 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_313_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_313_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_313 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_314_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_314_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_314 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_315_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_315_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_315 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_316_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_316_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_316 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_317_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_317_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_317 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_318_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_318_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_318 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_319_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_319_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_319 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_32_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_32_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_32 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_320_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_320_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_320 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_321_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_321_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_321 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_322_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_322_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_322 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_323_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_323_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_323 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_324_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_324_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_324 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_325_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_325_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_325 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_326_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_326_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_326 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_327_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_327_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_327 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_328_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_328_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_328 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_329_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_329_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_329 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_33_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_33_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_33 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_330_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_330_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_330 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_331_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_331_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_331 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_332_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_332_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_332 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_333_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_333_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_333 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_334_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_334_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_334 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_335_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_335_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_335 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_336_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_336_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_336 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_337_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_337_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_337 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_338_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_338_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_338 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_339_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_339_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_339 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_340_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_340_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_340 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_341_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_341_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_341 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_342_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_342_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_342 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_343_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_343_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_343 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_344_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_344_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_344 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_35_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_35_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_35 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_352_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_352_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_352 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_353_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_353_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_353 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_354_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_354_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_354 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_355_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_355_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_355 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_356_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_356_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_356 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_357_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_357_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_357 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_358_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_358_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_358 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_359_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_359_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_359 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_360_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_360_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_360 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_361_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_361_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_361 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_362_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_362_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_362 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_363_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_363_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_363 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_364_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_364_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_364 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_365_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_365_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_365 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_366_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_366_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_366 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_367_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_367_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_367 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_368_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_368_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_368 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_369_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_369_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_369 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_37_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_37_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_37 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_370_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_370_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_370 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_371_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_371_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_371 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_372_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_372_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_372 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_373_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_373_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_373 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_374_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_374_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_374 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_375_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_375_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_375 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_376_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_376_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_376 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_377_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_377_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_377 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_378_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_378_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_378 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_379_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_379_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_379 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_38_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_38_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_38 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_380_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_380_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_380 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_381_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_381_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_381 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_382_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_382_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_382 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_383_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_383_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_383 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_384_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_384_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_384 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_385_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_385_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_385 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_386_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_386_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_386 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_387_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_387_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_387 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_388_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_388_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_388 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_389_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_389_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_389 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_39_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_39_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_39 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_390_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_390_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_390 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_391_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_391_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_391 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_392_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_392_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_392 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_393_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_393_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_393 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_407_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_407_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_407 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_408_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_408_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_408 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_409_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_409_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_409 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_41_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_41_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_41 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_410_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_410_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_410 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_411_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_411_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_411 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_412_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_412_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_412 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_43_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_43_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_43 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_436_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_436_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_436 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_437_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_437_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_437 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_438_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_438_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_438 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_45_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_45_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_45 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_47_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_47_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_47 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_49_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_49_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_49 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_5_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_5_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_5 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_51_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_51_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_51 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_53_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_53_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_53 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_537_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_537_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_537 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_538_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_538_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_538 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_539_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_539_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_539 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_540_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_540_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_540 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_55_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_55_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_55 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_57_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_57_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_57 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_583_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_583_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_583 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_584_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_584_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_584 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_585_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_585_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_585 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_586_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_586_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_586 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_587_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_587_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_587 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_588_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_588_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_588 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_589_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_589_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_589 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_59_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_59_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_59 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_593_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_593_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_593 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_594_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_594_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_594 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_595_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_595_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_595 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_596_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_596_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_596 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_597_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_597_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_597 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_598_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_598_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_598 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_599_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_599_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_599 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_600_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_600_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_600 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_601_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_601_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_601 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_602_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_602_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_602 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_603_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_603_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_603 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_604_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_604_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_604 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_605_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_605_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_605 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_606_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_606_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_606 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_607_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_607_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_607 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_608_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_608_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_608 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_609_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_609_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_609 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_61_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_61_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_61 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_610_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_610_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_610 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_611_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_611_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_611 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_612_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_612_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_612 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_613_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_613_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_613 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_614_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_614_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_614 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_615_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_615_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_615 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_616_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_616_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_616 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_617_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_617_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_617 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_618_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_618_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_618 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_619_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_619_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_619 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_620_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_620_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_620 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_621_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_621_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_621 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_622_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_622_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_622 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_623_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_623_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_623 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_624_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_624_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_624 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_625_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_625_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_625 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_626_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_626_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_626 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_627_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_627_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_627 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_628_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_628_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_628 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_629_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_629_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_629 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_63_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_63_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_63 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_630_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_630_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_630 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_631_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_631_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_631 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_632_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_632_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_632 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_633_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_633_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_633 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_634_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_634_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_634 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_635_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_635_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_635 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_636_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_636_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_636 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_637_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_637_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_637 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_638_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_638_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_638 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_65_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_65_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_65 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_67_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_67_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_67 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_69_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_69_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_69 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_7_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_7_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_7 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_71_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_71_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_71 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_73_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_73_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_73 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_75_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_75_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_75 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_77_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_77_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_77 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_79_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_79_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_79 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_81_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_81_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_81 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_83_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_83_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_83 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_85_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_85_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_85 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_87_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_87_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_87 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_89_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_89_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_89 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_9_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_9_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_9 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_91_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_91_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_91 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_93_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_93_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_93 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_95_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_95_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_95 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_97_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_97_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_97 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_99_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._csignals_T_99_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._csignals_T_99 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_11_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_11_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_11 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_13_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_13_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_13 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_15_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_15_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_15 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_18_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_18_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_18 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_19_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_19_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_19 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_20_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_20_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_20 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_21_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_21_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_21 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_22_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_22_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_22 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_23_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_23_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_23 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_24_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_24_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_24 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_25_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_25_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_25 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_26_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_26_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_26 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_3_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_3_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_3 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_5_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_5_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_5 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_8_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_8_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._ctrl_pc_sel_no_xept_T_8 ;
	assign \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T ;
	assign \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_1_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_1 ;
	assign \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_2_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_2_obs_trg_arg0 = \Core_2stage.CtlPath_2stage._io_ctl_exception_cause_T_2 ;
	assign \Core_2stage.CtlPath_2stage.cs0_0_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.cs0_0_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.cs0_0 ;
	assign \Core_2stage.CtlPath_2stage.cs0_1_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.cs0_1_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.cs0_1 ;
	assign \Core_2stage.CtlPath_2stage.cs0_2_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.cs0_2_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.cs0_2 ;
	assign \Core_2stage.CtlPath_2stage.cs0_4_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.cs0_4_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.cs0_4 ;
	assign \Core_2stage.CtlPath_2stage.cs_alu_fun_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.cs_alu_fun_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.cs_alu_fun ;
	assign \Core_2stage.CtlPath_2stage.cs_br_type_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.cs_br_type_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.cs_br_type ;
	assign \Core_2stage.CtlPath_2stage.cs_val_inst_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.cs_val_inst_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.cs_val_inst ;
	assign \Core_2stage.CtlPath_2stage.csr_cmd_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.csr_cmd_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.csr_cmd ;
	assign \Core_2stage.CtlPath_2stage.csr_ren_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.csr_ren_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.csr_ren ;
	assign \Core_2stage.CtlPath_2stage.ctrl_pc_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.ctrl_pc_sel_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.ctrl_pc_sel ;
	assign \Core_2stage.CtlPath_2stage.ctrl_pc_sel_no_xept_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.ctrl_pc_sel_no_xept_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.ctrl_pc_sel_no_xept ;
	assign \Core_2stage.CtlPath_2stage.illegal_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.illegal_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.illegal ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_alu_fun_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_alu_fun_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_ctl_alu_fun ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_csr_cmd_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_csr_cmd_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_ctl_csr_cmd ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_exception_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_exception_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_ctl_exception ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_exception_cause_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_exception_cause_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_ctl_exception_cause ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_if_kill_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_if_kill_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_ctl_if_kill ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_mem_fcn_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_mem_fcn_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_ctl_mem_fcn ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_mem_typ_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_mem_typ_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_ctl_mem_typ ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_mem_val_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_mem_val_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_ctl_mem_val ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_op1_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_op1_sel_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_ctl_op1_sel ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_op2_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_op2_sel_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_ctl_op2_sel ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_pc_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_pc_sel_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_ctl_pc_sel ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_pc_sel_no_xept_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_pc_sel_no_xept_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_ctl_pc_sel_no_xept ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_rf_wen_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_rf_wen_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_ctl_rf_wen ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_stall_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_stall_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_ctl_stall ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_wb_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_ctl_wb_sel_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_ctl_wb_sel ;
	assign \Core_2stage.CtlPath_2stage.io_dat_br_eq_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_dat_br_eq_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_dat_br_eq ;
	assign \Core_2stage.CtlPath_2stage.io_dat_br_lt_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_dat_br_lt_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_dat_br_lt ;
	assign \Core_2stage.CtlPath_2stage.io_dat_br_ltu_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_dat_br_ltu_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_dat_br_ltu ;
	assign \Core_2stage.CtlPath_2stage.io_dat_csr_eret_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_dat_csr_eret_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_dat_csr_eret ;
	assign \Core_2stage.CtlPath_2stage.io_dat_csr_interrupt_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_dat_csr_interrupt_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_dat_csr_interrupt ;
	assign \Core_2stage.CtlPath_2stage.io_dat_data_misaligned_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_dat_data_misaligned_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_dat_data_misaligned ;
	assign \Core_2stage.CtlPath_2stage.io_dat_if_valid_resp_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_dat_if_valid_resp_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_dat_if_valid_resp ;
	assign \Core_2stage.CtlPath_2stage.io_dat_inst_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_dat_inst_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_dat_inst ;
	assign \Core_2stage.CtlPath_2stage.io_dat_inst_misaligned_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_dat_inst_misaligned_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_dat_inst_misaligned ;
	assign \Core_2stage.CtlPath_2stage.io_dat_mem_store_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_dat_mem_store_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_dat_mem_store ;
	assign \Core_2stage.CtlPath_2stage.io_dmem_req_bits_fcn_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_dmem_req_bits_fcn_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_dmem_req_bits_fcn ;
	assign \Core_2stage.CtlPath_2stage.io_dmem_req_bits_typ_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_dmem_req_bits_typ_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_dmem_req_bits_typ ;
	assign \Core_2stage.CtlPath_2stage.io_dmem_req_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_dmem_req_valid_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_dmem_req_valid ;
	assign \Core_2stage.CtlPath_2stage.io_dmem_resp_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_dmem_resp_valid_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_dmem_resp_valid ;
	assign \Core_2stage.CtlPath_2stage.io_imem_resp_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.io_imem_resp_valid_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.io_imem_resp_valid ;
	assign \Core_2stage.CtlPath_2stage.rs1_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.rs1_addr_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.rs1_addr ;
	assign \Core_2stage.CtlPath_2stage.stall_obs_trg_cond = 1 ;
	assign \Core_2stage.CtlPath_2stage.stall_obs_trg_arg0 = \Core_2stage.CtlPath_2stage.stall ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_0_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_0_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_0 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_145_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_145_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_145 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_146_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_146_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_146 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_170_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_170_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_170 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_174_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_174_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_174 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_175_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_175_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_175 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_176_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_176_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_176 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_178_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_178_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_178 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_180_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_180_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_180 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_182_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_182_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_182 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_183_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_183_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_183 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_2 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_207_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_207_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_207 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_211_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_211_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_211 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_212_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_212_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_212 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_213_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_213_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_213 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_215_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_215_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_215 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_217_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_217_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_217 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_239_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_239_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_239 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_241_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_241_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_241 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_242_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_242_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_242 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_273_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_273_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_273 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_274_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_274_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_274 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_279_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_279_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_279 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_293_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_293_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_293 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_294_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_294_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_294 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_296_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_296_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_296 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_298_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_298_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_298 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_3_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_3_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_3 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_300_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_300_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_300 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_315_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_315_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_315 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_316_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_316_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_316 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_318_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_318_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_318 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_34_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_34_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_34 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_341_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_341_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_341 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_342_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_342_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_342 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_343_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_343_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_343 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_344_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_344_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_344 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_345_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_345_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_345 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_346_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_346_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_346 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_35_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_35_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_35 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_40_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_40_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_40 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_41_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_41_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_41 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_46_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_46_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_46 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_48_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_48_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_48 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_51_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_51_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_51 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_52_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_52_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_52 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_73_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_73_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._GEN_73 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_14_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_14_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_14 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_15_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_15_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_15 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1714_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1714_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1714 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1717_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1717_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1717 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1719_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1719_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1719 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_172_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_172_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_172 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1722_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1722_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_1722 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_173_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_173_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_173 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_174_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_174_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_174 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_176_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_176_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_176 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_177_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_177_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_177 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_179_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_179_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_179 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_18_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_18_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_18 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_180_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_180_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_180 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_182_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_182_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_182 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_183_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_183_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_183 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_185_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_185_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_185 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_186_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_186_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_186 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_21_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_21_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_21 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_214_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_214_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_214 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_216_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_216_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_216 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_218_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_218_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_218 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_22_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_22_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_22 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_222_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_222_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_222 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_23_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_23_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_23 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_24_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_24_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_24 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_27_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_27_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_27 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_28_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_28_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_28 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_366_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_366_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_366 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_367_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_367_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_367 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_368_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._T_368_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._T_368 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._any_T_78_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._any_T_78_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._any_T_78 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugBreak_T_3_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugBreak_T_3_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugBreak_T_3 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugBreak_T_4_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugBreak_T_4_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugBreak_T_4 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugInt_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugInt_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugInt_T_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugTrigger_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugTrigger_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._causeIsDebugTrigger_T_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._cause_T_5_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._cause_T_5_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._cause_T_5 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._debugTVec_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._debugTVec_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._debugTVec_T ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_12_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_12_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_12 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_122_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_122_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_122 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_14_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_14_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_14 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_18_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_18_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_18 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_20_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_20_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_20 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_214_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_214_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_214 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_22_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_22_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_22 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_26_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_26_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_26 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_28_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_28_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_28 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_30_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_30_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_30 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_32_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_32_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_32 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_34_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_34_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_34 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_36_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_36_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_36 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_38_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_38_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_38 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_8_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_8_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._decoded_T_8 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._epc_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._epc_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._epc_T ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._epc_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._epc_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._epc_T_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_decode_0_read_illegal_T_16_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_decode_0_read_illegal_T_16_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_decode_0_read_illegal_T_16 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_eret_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_eret_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_eret_T ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_interrupt_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_interrupt_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_interrupt_T ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_10_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_10_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_10 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_107_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_107_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_107 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_108_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_108_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_108 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_11_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_11_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_11 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_115_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_115_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_115 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_116_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_116_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_116 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_117_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_117_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_117 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_118_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_118_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_118 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_119_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_119_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_119 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_12_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_12_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_12 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_120_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_120_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_120 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_121_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_121_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_121 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_122_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_122_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_122 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_123_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_123_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_123 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_124_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_124_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_124 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_125_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_125_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_125 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_126_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_126_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_126 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_127_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_127_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_127 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_128_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_128_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_128 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_129_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_129_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_129 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_13_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_13_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_13 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_130_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_130_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_130 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_14_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_14_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_14 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_15_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_15_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_15 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_16_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_16_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_16 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_17_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_17_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_17 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_18_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_18_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_18 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_19_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_19_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_19 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_218_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_218_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_218 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_219_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_219_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_219 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_4_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_4_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_4 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_5_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_5_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_5 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_6_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_6_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_6 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_7_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_7_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_7 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_8_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_8_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_8 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_9_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_9_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._io_rw_rdata_T_9 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._large_r_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._large_r_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._large_r_T_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._large_r_T_3_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._large_r_T_3_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._large_r_T_3 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._m_interrupts_T_3_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._m_interrupts_T_3_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._m_interrupts_T_3 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._m_interrupts_T_5_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._m_interrupts_T_5_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._m_interrupts_T_5 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._new_mstatus_WIRE_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._new_mstatus_WIRE_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._new_mstatus_WIRE ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._notDebugTVec_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._notDebugTVec_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._notDebugTVec_T_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mip_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mip_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mip_T ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mstatus_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mstatus_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mstatus_T ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_3_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_3_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_3 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_4_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_4_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._read_mtvec_T_4 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_dcsr_cause_T_2 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mcause_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mcause_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mcause_T ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mcountinhibit_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mcountinhibit_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mcountinhibit_T_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mepc_T_2 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mie_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mie_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._reg_mie_T ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_2 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_5_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_5_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_5 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_6_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_6_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._wdata_T_6 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_100_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_100_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_100 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_101_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_101_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_101 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_102_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_102_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_102 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_103_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_103_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_103 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_104_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_104_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_104 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_105_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_105_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_105 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_106_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_106_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_106 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_107_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_107_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_107 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_108_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_108_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_108 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_109_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_109_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_109 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_111_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_111_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_111 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_112_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_112_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_112 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_113_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_113_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_113 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_114_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_114_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_114 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_115_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_115_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_115 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_116_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_116_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_116 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_117_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_117_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_117 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_118_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_118_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_118 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_119_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_119_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_119 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_120_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_120_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_120 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_121_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_121_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_121 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_122_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_122_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_122 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_123_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_123_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_123 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_124_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_124_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_124 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_95_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_95_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_95 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_96_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_96_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_96 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_97_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_97_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_97 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_98_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_98_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_98 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_99_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_99_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage._which_T_99 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.addr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.addr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.addr ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.anyInterrupt_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.anyInterrupt_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.anyInterrupt ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.cause_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.cause_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.cause ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugBreak_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugBreak_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugBreak ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugInt_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugInt_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugInt ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugTrigger_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugTrigger_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.causeIsDebugTrigger ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.cause_lsbs_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.cause_lsbs_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.cause_lsbs ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.clock_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.clock_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.clock ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.csr_wen_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.csr_wen_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.csr_wen ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.d_interrupts_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.d_interrupts_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.d_interrupts ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.debugTVec_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.debugTVec_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.debugTVec ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_10_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_10_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_10 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_107_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_107_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_107 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_108_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_108_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_108 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_11_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_11_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_11 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_12_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_12_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_12 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_13_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_13_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_13 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_14_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_14_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_14 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_15_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_15_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_15 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_16_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_16_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_16 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_17_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_17_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_17 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_18_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_18_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_18 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_19_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_19_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_19 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_4_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_4_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_4 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_5_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_5_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_5 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_6_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_6_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_6 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_7_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_7_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_7 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_8_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_8_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_8 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_9_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_9_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.decoded_9 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.epc_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.epc_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.epc ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.exception_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.exception_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.exception ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_break_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_break_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_break ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_call_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_call_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_call ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_cease_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_cease_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_cease ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_ret_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_ret_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_ret ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_wfi_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_wfi_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.insn_wfi ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_cause_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_cause_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_cause ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_csr_stall_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_csr_stall_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_csr_stall ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_eret_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_eret_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_eret ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_evec_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_evec_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_evec ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_exception_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_exception_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_exception ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_hartid_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_hartid_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_hartid ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupt_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupt_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupt ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupt_cause_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupt_cause_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupt_cause ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_debug_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_debug_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_debug ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_meip_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_meip_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_meip ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_msip_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_msip_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_msip ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_mtip_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_mtip_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupts_mtip ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_pc_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_pc_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_pc ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_retire_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_retire_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_retire ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_addr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_addr ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_cmd_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_cmd_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_cmd ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_rdata_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_rdata_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_rdata ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_wdata_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_wdata_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_rw_wdata ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_singleStep_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_singleStep_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_singleStep ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease_r_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease_r_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease_r ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_debug_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_debug_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_debug ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_dprv_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_dprv_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_dprv ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_dv_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_dv_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_dv ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_fs_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_fs_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_fs ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_gva_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_gva_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_gva ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_hie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_hie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_hie ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_isa_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_isa_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_isa ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mbe_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mbe_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mbe ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mie ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpie ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpp_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpp_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpp ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mprv_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mprv_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mprv ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpv_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpv_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mpv ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mxr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mxr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_mxr ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_prv_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_prv_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_prv ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sbe_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sbe_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sbe ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sd_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sd_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sd ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sd_rv32_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sd_rv32_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sd_rv32 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sie ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_spie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_spie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_spie ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_spp_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_spp_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_spp ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sum_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sum_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sum ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sxl_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sxl_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_sxl ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tsr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tsr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tsr ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tvm_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tvm_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tvm ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tw_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tw_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_tw ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_ube_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_ube_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_ube ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_uie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_uie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_uie ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_upie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_upie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_upie ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_uxl_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_uxl_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_uxl ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_v_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_v_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_v ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_vs_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_vs_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_vs ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_wfi_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_wfi_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_wfi ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_xs_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_xs_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_xs ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_zero1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_zero1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_zero1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_zero2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_zero2_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_zero2 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_time_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_time_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_time ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_tval_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_tval_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_tval ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_ungated_clock_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_ungated_clock_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_ungated_clock ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.large__obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.large__obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.large_ ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.large_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.large_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.large_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.m_interrupts_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.m_interrupts_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.m_interrupts ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.new_dcsr_ebreakm_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.new_dcsr_ebreakm_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.new_dcsr_ebreakm ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.new_mstatus_mie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.new_mstatus_mie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.new_mstatus_mie ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.new_mstatus_mpie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.new_mstatus_mpie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.new_mstatus_mpie ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.nextSmall_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.nextSmall_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.nextSmall ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.nextSmall_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.nextSmall_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.nextSmall_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_doVector_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_doVector_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_doVector ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_interruptOffset_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_interruptOffset_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_interruptOffset ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_interruptVec_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_interruptVec_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.notDebugTVec_interruptVec ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.pending_interrupts_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.pending_interrupts_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.pending_interrupts ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mip_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mip_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mip ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_hi_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_hi_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_hi ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_hi_hi_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_hi_hi_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_hi_hi ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_lo_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_lo_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_lo ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_lo_lo_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_lo_lo_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mstatus_lo_lo ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mtvec_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mtvec_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.read_mtvec ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_cause_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_cause_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_cause ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_ebreakm_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_ebreakm_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_ebreakm ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_step_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_step_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_step ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_debug_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_debug_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_debug ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dpc_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dpc_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dpc ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dscratch_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dscratch_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dscratch ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcause_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcause_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcause ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcountinhibit_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcountinhibit_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcountinhibit ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mepc_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mepc_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mepc ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mie ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mscratch_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mscratch_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mscratch ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mie ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mpie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mpie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mpie ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_spp_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_spp_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_spp ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtval_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtval_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtval ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtvec_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtvec_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtvec ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_singleStepped_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_singleStepped_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_singleStepped ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_wfi_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_wfi_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_wfi ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reset_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reset_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.reset ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.small__obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.small__obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.small_ ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.small_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.small_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.small_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.system_insn_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.system_insn_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.system_insn ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.trapToDebug_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.trapToDebug_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.trapToDebug ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.tvec_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.tvec_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.tvec ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.value_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.value_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.value ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.value_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.value_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.value_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.wdata_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.wdata_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.wdata ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.whichInterrupt_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.whichInterrupt_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.whichInterrupt ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.x79_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.x79_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.x79 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.x86_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.x86_obs_trg_arg0 = \Core_2stage.DatPath_2stage.CSRFile_2stage.x86 ;
	assign \Core_2stage.DatPath_2stage._GEN_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._GEN_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage._GEN_1 ;
	assign \Core_2stage.DatPath_2stage._GEN_11_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._GEN_11_obs_trg_arg0 = \Core_2stage.DatPath_2stage._GEN_11 ;
	assign \Core_2stage.DatPath_2stage._GEN_3_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._GEN_3_obs_trg_arg0 = \Core_2stage.DatPath_2stage._GEN_3 ;
	assign \Core_2stage.DatPath_2stage._T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._T_obs_trg_arg0 = \Core_2stage.DatPath_2stage._T ;
	assign \Core_2stage.DatPath_2stage._T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage._T_1 ;
	assign \Core_2stage.DatPath_2stage._T_10_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._T_10_obs_trg_arg0 = \Core_2stage.DatPath_2stage._T_10 ;
	assign \Core_2stage.DatPath_2stage._T_12_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._T_12_obs_trg_arg0 = \Core_2stage.DatPath_2stage._T_12 ;
	assign \Core_2stage.DatPath_2stage._T_14_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._T_14_obs_trg_arg0 = \Core_2stage.DatPath_2stage._T_14 ;
	assign \Core_2stage.DatPath_2stage._T_16_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._T_16_obs_trg_arg0 = \Core_2stage.DatPath_2stage._T_16 ;
	assign \Core_2stage.DatPath_2stage._T_17_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._T_17_obs_trg_arg0 = \Core_2stage.DatPath_2stage._T_17 ;
	assign \Core_2stage.DatPath_2stage._T_4_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._T_4_obs_trg_arg0 = \Core_2stage.DatPath_2stage._T_4 ;
	assign \Core_2stage.DatPath_2stage._T_5_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._T_5_obs_trg_arg0 = \Core_2stage.DatPath_2stage._T_5 ;
	assign \Core_2stage.DatPath_2stage._T_6_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._T_6_obs_trg_arg0 = \Core_2stage.DatPath_2stage._T_6 ;
	assign \Core_2stage.DatPath_2stage._T_8_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._T_8_obs_trg_arg0 = \Core_2stage.DatPath_2stage._T_8 ;
	assign \Core_2stage.DatPath_2stage._csr_io_tval_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._csr_io_tval_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage._csr_io_tval_T ;
	assign \Core_2stage.DatPath_2stage._csr_io_tval_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._csr_io_tval_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage._csr_io_tval_T_1 ;
	assign \Core_2stage.DatPath_2stage._csr_io_tval_T_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._csr_io_tval_T_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage._csr_io_tval_T_2 ;
	assign \Core_2stage.DatPath_2stage._csr_io_tval_T_3_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._csr_io_tval_T_3_obs_trg_arg0 = \Core_2stage.DatPath_2stage._csr_io_tval_T_3 ;
	assign \Core_2stage.DatPath_2stage._csr_io_tval_T_4_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._csr_io_tval_T_4_obs_trg_arg0 = \Core_2stage.DatPath_2stage._csr_io_tval_T_4 ;
	assign \Core_2stage.DatPath_2stage._csr_io_tval_T_5_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._csr_io_tval_T_5_obs_trg_arg0 = \Core_2stage.DatPath_2stage._csr_io_tval_T_5 ;
	assign \Core_2stage.DatPath_2stage._csr_io_tval_T_6_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._csr_io_tval_T_6_obs_trg_arg0 = \Core_2stage.DatPath_2stage._csr_io_tval_T_6 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op1_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op1_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_op1_T ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op1_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op1_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_op1_T_1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op1_T_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op1_T_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_op1_T_2 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op1_T_3_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op1_T_3_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_op1_T_3 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op1_T_4_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op1_T_4_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_op1_T_4 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op2_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op2_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_op2_T ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op2_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op2_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_op2_T_1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op2_T_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op2_T_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_op2_T_2 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op2_T_3_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op2_T_3_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_op2_T_3 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op2_T_4_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op2_T_4_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_op2_T_4 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op2_T_5_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op2_T_5_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_op2_T_5 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op2_T_6_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_op2_T_6_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_op2_T_6 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_10_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_10_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_10 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_11_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_11_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_11 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_12_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_12_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_12 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_13_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_13_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_13 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_14_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_14_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_14 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_15_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_15_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_15 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_16_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_16_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_16 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_17_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_17_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_17 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_18_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_18_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_18 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_19_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_19_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_19 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_2 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_21_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_21_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_21 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_24_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_24_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_24 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_25_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_25_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_25 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_26_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_26_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_26 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_27_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_27_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_27 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_28_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_28_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_28 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_29_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_29_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_29 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_3_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_3_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_3 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_30_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_30_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_30 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_31_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_31_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_31 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_32_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_32_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_32 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_33_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_33_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_33 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_34_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_34_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_34 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_35_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_35_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_35 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_36_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_36_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_36 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_37_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_37_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_37 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_5_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_5_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_5 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_6_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_6_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_6 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_7_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_7_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_7 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_8_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_8_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_8 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_9_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_alu_out_T_9_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_alu_out_T_9 ;
	assign \Core_2stage.DatPath_2stage._exe_jump_reg_target_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_jump_reg_target_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_jump_reg_target_T_1 ;
	assign \Core_2stage.DatPath_2stage._exe_wbdata_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_wbdata_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_wbdata_T ;
	assign \Core_2stage.DatPath_2stage._exe_wbdata_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_wbdata_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_wbdata_T_1 ;
	assign \Core_2stage.DatPath_2stage._exe_wbdata_T_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_wbdata_T_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_wbdata_T_2 ;
	assign \Core_2stage.DatPath_2stage._exe_wbdata_T_3_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_wbdata_T_3_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_wbdata_T_3 ;
	assign \Core_2stage.DatPath_2stage._exe_wbdata_T_4_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_wbdata_T_4_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_wbdata_T_4 ;
	assign \Core_2stage.DatPath_2stage._exe_wbdata_T_5_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_wbdata_T_5_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_wbdata_T_5 ;
	assign \Core_2stage.DatPath_2stage._exe_wbdata_T_6_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._exe_wbdata_T_6_obs_trg_arg0 = \Core_2stage.DatPath_2stage._exe_wbdata_T_6 ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage._if_pc_next_T ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage._if_pc_next_T_1 ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage._if_pc_next_T_2 ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_3_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_3_obs_trg_arg0 = \Core_2stage.DatPath_2stage._if_pc_next_T_3 ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_4_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_4_obs_trg_arg0 = \Core_2stage.DatPath_2stage._if_pc_next_T_4 ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_5_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_5_obs_trg_arg0 = \Core_2stage.DatPath_2stage._if_pc_next_T_5 ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_6_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_6_obs_trg_arg0 = \Core_2stage.DatPath_2stage._if_pc_next_T_6 ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_7_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._if_pc_next_T_7_obs_trg_arg0 = \Core_2stage.DatPath_2stage._if_pc_next_T_7 ;
	assign \Core_2stage.DatPath_2stage._imm_b_sext_T_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._imm_b_sext_T_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage._imm_b_sext_T_2 ;
	assign \Core_2stage.DatPath_2stage._imm_i_sext_T_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._imm_i_sext_T_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage._imm_i_sext_T_2 ;
	assign \Core_2stage.DatPath_2stage._imm_j_sext_T_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._imm_j_sext_T_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage._imm_j_sext_T_2 ;
	assign \Core_2stage.DatPath_2stage._imm_s_sext_T_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._imm_s_sext_T_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage._imm_s_sext_T_2 ;
	assign \Core_2stage.DatPath_2stage._io_dat_br_lt_T_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._io_dat_br_lt_T_obs_trg_arg0 = \Core_2stage.DatPath_2stage._io_dat_br_lt_T ;
	assign \Core_2stage.DatPath_2stage._io_dat_br_lt_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._io_dat_br_lt_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage._io_dat_br_lt_T_1 ;
	assign \Core_2stage.DatPath_2stage._io_dat_data_misaligned_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._io_dat_data_misaligned_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage._io_dat_data_misaligned_T_1 ;
	assign \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_11_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_11_obs_trg_arg0 = \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_11 ;
	assign \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_12_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_12_obs_trg_arg0 = \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_12 ;
	assign \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_2_obs_trg_arg0 = \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_2 ;
	assign \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_6_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_6_obs_trg_arg0 = \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_6 ;
	assign \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_7_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_7_obs_trg_arg0 = \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_7 ;
	assign \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_8_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_8_obs_trg_arg0 = \Core_2stage.DatPath_2stage._io_dat_inst_misaligned_T_8 ;
	assign \Core_2stage.DatPath_2stage._misaligned_mask_T_1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._misaligned_mask_T_1_obs_trg_arg0 = \Core_2stage.DatPath_2stage._misaligned_mask_T_1 ;
	assign \Core_2stage.DatPath_2stage._misaligned_mask_T_3_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._misaligned_mask_T_3_obs_trg_arg0 = \Core_2stage.DatPath_2stage._misaligned_mask_T_3 ;
	assign \Core_2stage.DatPath_2stage._misaligned_mask_T_4_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._misaligned_mask_T_4_obs_trg_arg0 = \Core_2stage.DatPath_2stage._misaligned_mask_T_4 ;
	assign \Core_2stage.DatPath_2stage._tval_inst_ma_T_3_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._tval_inst_ma_T_3_obs_trg_arg0 = \Core_2stage.DatPath_2stage._tval_inst_ma_T_3 ;
	assign \Core_2stage.DatPath_2stage._tval_inst_ma_T_4_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage._tval_inst_ma_T_4_obs_trg_arg0 = \Core_2stage.DatPath_2stage._tval_inst_ma_T_4 ;
	assign \Core_2stage.DatPath_2stage.alu_shamt_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.alu_shamt_obs_trg_arg0 = \Core_2stage.DatPath_2stage.alu_shamt ;
	assign \Core_2stage.DatPath_2stage.clock_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.clock_obs_trg_arg0 = \Core_2stage.DatPath_2stage.clock ;
	assign \Core_2stage.DatPath_2stage.csr_clock_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_clock_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_clock ;
	assign \Core_2stage.DatPath_2stage.csr_io_cause_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_cause_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_cause ;
	assign \Core_2stage.DatPath_2stage.csr_io_csr_stall_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_csr_stall_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_csr_stall ;
	assign \Core_2stage.DatPath_2stage.csr_io_eret_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_eret_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_eret ;
	assign \Core_2stage.DatPath_2stage.csr_io_evec_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_evec_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_evec ;
	assign \Core_2stage.DatPath_2stage.csr_io_exception_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_exception_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_exception ;
	assign \Core_2stage.DatPath_2stage.csr_io_hartid_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_hartid_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_hartid ;
	assign \Core_2stage.DatPath_2stage.csr_io_interrupt_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_interrupt_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_interrupt ;
	assign \Core_2stage.DatPath_2stage.csr_io_interrupt_cause_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_interrupt_cause_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_interrupt_cause ;
	assign \Core_2stage.DatPath_2stage.csr_io_interrupts_debug_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_interrupts_debug_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_interrupts_debug ;
	assign \Core_2stage.DatPath_2stage.csr_io_interrupts_meip_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_interrupts_meip_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_interrupts_meip ;
	assign \Core_2stage.DatPath_2stage.csr_io_interrupts_msip_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_interrupts_msip_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_interrupts_msip ;
	assign \Core_2stage.DatPath_2stage.csr_io_interrupts_mtip_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_interrupts_mtip_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_interrupts_mtip ;
	assign \Core_2stage.DatPath_2stage.csr_io_pc_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_pc_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_pc ;
	assign \Core_2stage.DatPath_2stage.csr_io_retire_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_retire_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_retire ;
	assign \Core_2stage.DatPath_2stage.csr_io_rw_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_rw_addr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_rw_addr ;
	assign \Core_2stage.DatPath_2stage.csr_io_rw_cmd_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_rw_cmd_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_rw_cmd ;
	assign \Core_2stage.DatPath_2stage.csr_io_rw_rdata_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_rw_rdata_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_rw_rdata ;
	assign \Core_2stage.DatPath_2stage.csr_io_rw_wdata_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_rw_wdata_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_rw_wdata ;
	assign \Core_2stage.DatPath_2stage.csr_io_singleStep_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_singleStep_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_singleStep ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_cease_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_cease_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_cease ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_debug_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_debug_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_debug ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_dprv_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_dprv_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_dprv ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_dv_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_dv_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_dv ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_fs_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_fs_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_fs ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_gva_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_gva_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_gva ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_hie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_hie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_hie ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_isa_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_isa_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_isa ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_mbe_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_mbe_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_mbe ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_mie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_mie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_mie ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_mpie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_mpie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_mpie ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_mpp_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_mpp_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_mpp ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_mprv_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_mprv_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_mprv ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_mpv_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_mpv_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_mpv ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_mxr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_mxr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_mxr ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_prv_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_prv_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_prv ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_sbe_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_sbe_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_sbe ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_sd_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_sd_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_sd ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_sd_rv32_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_sd_rv32_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_sd_rv32 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_sie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_sie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_sie ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_spie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_spie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_spie ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_spp_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_spp_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_spp ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_sum_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_sum_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_sum ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_sxl_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_sxl_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_sxl ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_tsr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_tsr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_tsr ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_tvm_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_tvm_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_tvm ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_tw_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_tw_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_tw ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_ube_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_ube_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_ube ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_uie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_uie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_uie ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_upie_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_upie_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_upie ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_uxl_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_uxl_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_uxl ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_v_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_v_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_v ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_vs_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_vs_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_vs ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_wfi_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_wfi_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_wfi ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_xs_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_xs_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_xs ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_zero1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_zero1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_zero1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_zero2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_status_zero2_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_status_zero2 ;
	assign \Core_2stage.DatPath_2stage.csr_io_time_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_time_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_time ;
	assign \Core_2stage.DatPath_2stage.csr_io_tval_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_tval_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_tval ;
	assign \Core_2stage.DatPath_2stage.csr_io_ungated_clock_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_io_ungated_clock_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_io_ungated_clock ;
	assign \Core_2stage.DatPath_2stage.csr_reset_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.csr_reset_obs_trg_arg0 = \Core_2stage.DatPath_2stage.csr_reset ;
	assign \Core_2stage.DatPath_2stage.decode_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.decode_obs_trg_arg0 = \Core_2stage.DatPath_2stage.decode ;
	assign \Core_2stage.DatPath_2stage.exception_target_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exception_target_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exception_target ;
	assign \Core_2stage.DatPath_2stage.exe_alu_op1_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_alu_op1_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_alu_op1 ;
	assign \Core_2stage.DatPath_2stage.exe_alu_op2_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_alu_op2_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_alu_op2 ;
	assign \Core_2stage.DatPath_2stage.exe_alu_out_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_alu_out_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_alu_out ;
	assign \Core_2stage.DatPath_2stage.exe_br_target_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_br_target_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_br_target ;
	assign \Core_2stage.DatPath_2stage.exe_jmp_target_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_jmp_target_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_jmp_target ;
	assign \Core_2stage.DatPath_2stage.exe_jump_reg_target_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_jump_reg_target_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_jump_reg_target ;
	assign \Core_2stage.DatPath_2stage.exe_reg_inst_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_reg_inst_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_reg_inst ;
	assign \Core_2stage.DatPath_2stage.exe_reg_pc_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_reg_pc_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_reg_pc ;
	assign \Core_2stage.DatPath_2stage.exe_reg_pc_plus4_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_reg_pc_plus4_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_reg_pc_plus4 ;
	assign \Core_2stage.DatPath_2stage.exe_reg_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_reg_valid_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_reg_valid ;
	assign \Core_2stage.DatPath_2stage.exe_rs1_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_rs1_addr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_rs1_addr ;
	assign \Core_2stage.DatPath_2stage.exe_rs1_data_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_rs1_data_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_rs1_data ;
	assign \Core_2stage.DatPath_2stage.exe_rs2_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_rs2_addr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_rs2_addr ;
	assign \Core_2stage.DatPath_2stage.exe_rs2_data_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_rs2_data_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_rs2_data ;
	assign \Core_2stage.DatPath_2stage.exe_wbaddr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_wbaddr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_wbaddr ;
	assign \Core_2stage.DatPath_2stage.exe_wbdata_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_wbdata_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_wbdata ;
	assign \Core_2stage.DatPath_2stage.exe_wben_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.exe_wben_obs_trg_arg0 = \Core_2stage.DatPath_2stage.exe_wben ;
	assign \Core_2stage.DatPath_2stage.if_inst_buffer_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.if_inst_buffer_obs_trg_arg0 = \Core_2stage.DatPath_2stage.if_inst_buffer ;
	assign \Core_2stage.DatPath_2stage.if_inst_buffer_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.if_inst_buffer_valid_obs_trg_arg0 = \Core_2stage.DatPath_2stage.if_inst_buffer_valid ;
	assign \Core_2stage.DatPath_2stage.if_pc_plus4_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.if_pc_plus4_obs_trg_arg0 = \Core_2stage.DatPath_2stage.if_pc_plus4 ;
	assign \Core_2stage.DatPath_2stage.if_reg_pc_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.if_reg_pc_obs_trg_arg0 = \Core_2stage.DatPath_2stage.if_reg_pc ;
	assign \Core_2stage.DatPath_2stage.imm_b_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.imm_b_obs_trg_arg0 = \Core_2stage.DatPath_2stage.imm_b ;
	assign \Core_2stage.DatPath_2stage.imm_b_sext_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.imm_b_sext_obs_trg_arg0 = \Core_2stage.DatPath_2stage.imm_b_sext ;
	assign \Core_2stage.DatPath_2stage.imm_i_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.imm_i_obs_trg_arg0 = \Core_2stage.DatPath_2stage.imm_i ;
	assign \Core_2stage.DatPath_2stage.imm_i_sext_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.imm_i_sext_obs_trg_arg0 = \Core_2stage.DatPath_2stage.imm_i_sext ;
	assign \Core_2stage.DatPath_2stage.imm_j_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.imm_j_obs_trg_arg0 = \Core_2stage.DatPath_2stage.imm_j ;
	assign \Core_2stage.DatPath_2stage.imm_j_sext_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.imm_j_sext_obs_trg_arg0 = \Core_2stage.DatPath_2stage.imm_j_sext ;
	assign \Core_2stage.DatPath_2stage.imm_s_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.imm_s_obs_trg_arg0 = \Core_2stage.DatPath_2stage.imm_s ;
	assign \Core_2stage.DatPath_2stage.imm_s_sext_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.imm_s_sext_obs_trg_arg0 = \Core_2stage.DatPath_2stage.imm_s_sext ;
	assign \Core_2stage.DatPath_2stage.imm_u_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.imm_u_obs_trg_arg0 = \Core_2stage.DatPath_2stage.imm_u ;
	assign \Core_2stage.DatPath_2stage.imm_u_sext_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.imm_u_sext_obs_trg_arg0 = \Core_2stage.DatPath_2stage.imm_u_sext ;
	assign \Core_2stage.DatPath_2stage.imm_z_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.imm_z_obs_trg_arg0 = \Core_2stage.DatPath_2stage.imm_z ;
	assign \Core_2stage.DatPath_2stage.io_ctl_alu_fun_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_alu_fun_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_alu_fun ;
	assign \Core_2stage.DatPath_2stage.io_ctl_csr_cmd_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_csr_cmd_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_csr_cmd ;
	assign \Core_2stage.DatPath_2stage.io_ctl_exception_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_exception_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_exception ;
	assign \Core_2stage.DatPath_2stage.io_ctl_exception_cause_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_exception_cause_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_exception_cause ;
	assign \Core_2stage.DatPath_2stage.io_ctl_if_kill_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_if_kill_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_if_kill ;
	assign \Core_2stage.DatPath_2stage.io_ctl_if_kill_r_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_if_kill_r_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_if_kill_r ;
	assign \Core_2stage.DatPath_2stage.io_ctl_mem_fcn_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_mem_fcn_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_mem_fcn ;
	assign \Core_2stage.DatPath_2stage.io_ctl_mem_typ_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_mem_typ_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_mem_typ ;
	assign \Core_2stage.DatPath_2stage.io_ctl_mem_val_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_mem_val_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_mem_val ;
	assign \Core_2stage.DatPath_2stage.io_ctl_op1_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_op1_sel_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_op1_sel ;
	assign \Core_2stage.DatPath_2stage.io_ctl_op2_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_op2_sel_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_op2_sel ;
	assign \Core_2stage.DatPath_2stage.io_ctl_pc_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_pc_sel_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_pc_sel ;
	assign \Core_2stage.DatPath_2stage.io_ctl_pc_sel_no_xept_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_pc_sel_no_xept_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_pc_sel_no_xept ;
	assign \Core_2stage.DatPath_2stage.io_ctl_rf_wen_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_rf_wen_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_rf_wen ;
	assign \Core_2stage.DatPath_2stage.io_ctl_stall_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_stall_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_stall ;
	assign \Core_2stage.DatPath_2stage.io_ctl_wb_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_ctl_wb_sel_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_ctl_wb_sel ;
	assign \Core_2stage.DatPath_2stage.io_dat_br_eq_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_dat_br_eq_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_dat_br_eq ;
	assign \Core_2stage.DatPath_2stage.io_dat_br_lt_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_dat_br_lt_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_dat_br_lt ;
	assign \Core_2stage.DatPath_2stage.io_dat_br_ltu_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_dat_br_ltu_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_dat_br_ltu ;
	assign \Core_2stage.DatPath_2stage.io_dat_csr_eret_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_dat_csr_eret_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_dat_csr_eret ;
	assign \Core_2stage.DatPath_2stage.io_dat_csr_interrupt_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_dat_csr_interrupt_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_dat_csr_interrupt ;
	assign \Core_2stage.DatPath_2stage.io_dat_data_misaligned_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_dat_data_misaligned_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_dat_data_misaligned ;
	assign \Core_2stage.DatPath_2stage.io_dat_if_valid_resp_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_dat_if_valid_resp_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_dat_if_valid_resp ;
	assign \Core_2stage.DatPath_2stage.io_dat_inst_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_dat_inst_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_dat_inst ;
	assign \Core_2stage.DatPath_2stage.io_dat_inst_misaligned_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_dat_inst_misaligned_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_dat_inst_misaligned ;
	assign \Core_2stage.DatPath_2stage.io_dat_mem_store_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_dat_mem_store_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_dat_mem_store ;
	assign \Core_2stage.DatPath_2stage.io_dmem_req_bits_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_dmem_req_bits_addr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_dmem_req_bits_addr ;
	assign \Core_2stage.DatPath_2stage.io_dmem_req_bits_data_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_dmem_req_bits_data_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_dmem_req_bits_data ;
	assign \Core_2stage.DatPath_2stage.io_dmem_resp_bits_data_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_dmem_resp_bits_data_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_dmem_resp_bits_data ;
	assign \Core_2stage.DatPath_2stage.io_hartid_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_hartid_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_hartid ;
	assign \Core_2stage.DatPath_2stage.io_imem_req_bits_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_imem_req_bits_addr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_imem_req_bits_addr ;
	assign \Core_2stage.DatPath_2stage.io_imem_req_bits_addr_state_invariant_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_imem_req_bits_addr_state_invariant_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_imem_req_bits_addr_state_invariant ;
	assign \Core_2stage.DatPath_2stage.io_imem_req_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_imem_req_valid_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_imem_req_valid ;
	assign \Core_2stage.DatPath_2stage.io_imem_resp_bits_data_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_imem_resp_bits_data_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_imem_resp_bits_data ;
	assign \Core_2stage.DatPath_2stage.io_imem_resp_bits_data_state_invariant_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_imem_resp_bits_data_state_invariant_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_imem_resp_bits_data_state_invariant ;
	assign \Core_2stage.DatPath_2stage.io_imem_resp_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_imem_resp_valid_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_imem_resp_valid ;
	assign \Core_2stage.DatPath_2stage.io_interrupt_debug_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_interrupt_debug_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_interrupt_debug ;
	assign \Core_2stage.DatPath_2stage.io_interrupt_meip_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_interrupt_meip_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_interrupt_meip ;
	assign \Core_2stage.DatPath_2stage.io_interrupt_msip_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_interrupt_msip_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_interrupt_msip ;
	assign \Core_2stage.DatPath_2stage.io_interrupt_mtip_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_interrupt_mtip_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_interrupt_mtip ;
	assign \Core_2stage.DatPath_2stage.io_reset_vector_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.io_reset_vector_obs_trg_arg0 = \Core_2stage.DatPath_2stage.io_reset_vector ;
	assign \Core_2stage.DatPath_2stage.misaligned_mask_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.misaligned_mask_obs_trg_arg0 = \Core_2stage.DatPath_2stage.misaligned_mask ;
	assign \Core_2stage.DatPath_2stage.pc_x_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.pc_x_obs_trg_arg0 = \Core_2stage.DatPath_2stage.pc_x ;
	assign \Core_2stage.DatPath_2stage.reg_interrupt_handled_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.reg_interrupt_handled_obs_trg_arg0 = \Core_2stage.DatPath_2stage.reg_interrupt_handled ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_1_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_1_addr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_MPORT_1_addr ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_1_data_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_1_data_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_MPORT_1_data ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_1_en_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_1_en_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_MPORT_1_en ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_1_mask_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_1_mask_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_MPORT_1_mask ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_addr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_MPORT_addr ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_data_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_data_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_MPORT_data ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_en_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_en_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_MPORT_en ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_mask_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_MPORT_mask_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_MPORT_mask ;
	assign \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_addr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_addr ;
	assign \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_data_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_data_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_data ;
	assign \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_en_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_en_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_exe_rs1_data_MPORT_en ;
	assign \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_addr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_addr ;
	assign \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_data_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_data_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_data ;
	assign \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_en_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_en_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_exe_rs2_data_MPORT_en ;
	assign \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_addr_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_addr ;
	assign \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_data_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_data_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_data ;
	assign \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_en_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_en_obs_trg_arg0 = \Core_2stage.DatPath_2stage.regfile_io_ddpath_rdata_MPORT_en ;
	assign \Core_2stage.DatPath_2stage.reset_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.reset_obs_trg_arg0 = \Core_2stage.DatPath_2stage.reset ;
	assign \Core_2stage.DatPath_2stage.tval_inst_ma_obs_trg_cond = 1 ;
	assign \Core_2stage.DatPath_2stage.tval_inst_ma_obs_trg_arg0 = \Core_2stage.DatPath_2stage.tval_inst_ma ;
	assign \Core_2stage.c_io_ctl_alu_fun_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_ctl_alu_fun_obs_trg_arg0 = \Core_2stage.c_io_ctl_alu_fun ;
	assign \Core_2stage.c_io_ctl_csr_cmd_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_ctl_csr_cmd_obs_trg_arg0 = \Core_2stage.c_io_ctl_csr_cmd ;
	assign \Core_2stage.c_io_ctl_exception_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_ctl_exception_obs_trg_arg0 = \Core_2stage.c_io_ctl_exception ;
	assign \Core_2stage.c_io_ctl_exception_cause_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_ctl_exception_cause_obs_trg_arg0 = \Core_2stage.c_io_ctl_exception_cause ;
	assign \Core_2stage.c_io_ctl_if_kill_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_ctl_if_kill_obs_trg_arg0 = \Core_2stage.c_io_ctl_if_kill ;
	assign \Core_2stage.c_io_ctl_mem_fcn_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_ctl_mem_fcn_obs_trg_arg0 = \Core_2stage.c_io_ctl_mem_fcn ;
	assign \Core_2stage.c_io_ctl_mem_typ_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_ctl_mem_typ_obs_trg_arg0 = \Core_2stage.c_io_ctl_mem_typ ;
	assign \Core_2stage.c_io_ctl_mem_val_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_ctl_mem_val_obs_trg_arg0 = \Core_2stage.c_io_ctl_mem_val ;
	assign \Core_2stage.c_io_ctl_op1_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_ctl_op1_sel_obs_trg_arg0 = \Core_2stage.c_io_ctl_op1_sel ;
	assign \Core_2stage.c_io_ctl_op2_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_ctl_op2_sel_obs_trg_arg0 = \Core_2stage.c_io_ctl_op2_sel ;
	assign \Core_2stage.c_io_ctl_pc_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_ctl_pc_sel_obs_trg_arg0 = \Core_2stage.c_io_ctl_pc_sel ;
	assign \Core_2stage.c_io_ctl_pc_sel_no_xept_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_ctl_pc_sel_no_xept_obs_trg_arg0 = \Core_2stage.c_io_ctl_pc_sel_no_xept ;
	assign \Core_2stage.c_io_ctl_rf_wen_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_ctl_rf_wen_obs_trg_arg0 = \Core_2stage.c_io_ctl_rf_wen ;
	assign \Core_2stage.c_io_ctl_stall_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_ctl_stall_obs_trg_arg0 = \Core_2stage.c_io_ctl_stall ;
	assign \Core_2stage.c_io_ctl_wb_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_ctl_wb_sel_obs_trg_arg0 = \Core_2stage.c_io_ctl_wb_sel ;
	assign \Core_2stage.c_io_dat_br_eq_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_dat_br_eq_obs_trg_arg0 = \Core_2stage.c_io_dat_br_eq ;
	assign \Core_2stage.c_io_dat_br_lt_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_dat_br_lt_obs_trg_arg0 = \Core_2stage.c_io_dat_br_lt ;
	assign \Core_2stage.c_io_dat_br_ltu_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_dat_br_ltu_obs_trg_arg0 = \Core_2stage.c_io_dat_br_ltu ;
	assign \Core_2stage.c_io_dat_csr_eret_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_dat_csr_eret_obs_trg_arg0 = \Core_2stage.c_io_dat_csr_eret ;
	assign \Core_2stage.c_io_dat_csr_interrupt_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_dat_csr_interrupt_obs_trg_arg0 = \Core_2stage.c_io_dat_csr_interrupt ;
	assign \Core_2stage.c_io_dat_data_misaligned_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_dat_data_misaligned_obs_trg_arg0 = \Core_2stage.c_io_dat_data_misaligned ;
	assign \Core_2stage.c_io_dat_if_valid_resp_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_dat_if_valid_resp_obs_trg_arg0 = \Core_2stage.c_io_dat_if_valid_resp ;
	assign \Core_2stage.c_io_dat_inst_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_dat_inst_obs_trg_arg0 = \Core_2stage.c_io_dat_inst ;
	assign \Core_2stage.c_io_dat_inst_misaligned_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_dat_inst_misaligned_obs_trg_arg0 = \Core_2stage.c_io_dat_inst_misaligned ;
	assign \Core_2stage.c_io_dat_mem_store_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_dat_mem_store_obs_trg_arg0 = \Core_2stage.c_io_dat_mem_store ;
	assign \Core_2stage.c_io_dmem_req_bits_fcn_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_dmem_req_bits_fcn_obs_trg_arg0 = \Core_2stage.c_io_dmem_req_bits_fcn ;
	assign \Core_2stage.c_io_dmem_req_bits_typ_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_dmem_req_bits_typ_obs_trg_arg0 = \Core_2stage.c_io_dmem_req_bits_typ ;
	assign \Core_2stage.c_io_dmem_req_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_dmem_req_valid_obs_trg_arg0 = \Core_2stage.c_io_dmem_req_valid ;
	assign \Core_2stage.c_io_dmem_resp_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_dmem_resp_valid_obs_trg_arg0 = \Core_2stage.c_io_dmem_resp_valid ;
	assign \Core_2stage.c_io_imem_resp_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.c_io_imem_resp_valid_obs_trg_arg0 = \Core_2stage.c_io_imem_resp_valid ;
	assign \Core_2stage.clock_obs_trg_cond = 1 ;
	assign \Core_2stage.clock_obs_trg_arg0 = \Core_2stage.clock ;
	assign \Core_2stage.d_clock_obs_trg_cond = 1 ;
	assign \Core_2stage.d_clock_obs_trg_arg0 = \Core_2stage.d_clock ;
	assign \Core_2stage.d_io_ctl_alu_fun_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_ctl_alu_fun_obs_trg_arg0 = \Core_2stage.d_io_ctl_alu_fun ;
	assign \Core_2stage.d_io_ctl_csr_cmd_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_ctl_csr_cmd_obs_trg_arg0 = \Core_2stage.d_io_ctl_csr_cmd ;
	assign \Core_2stage.d_io_ctl_exception_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_ctl_exception_obs_trg_arg0 = \Core_2stage.d_io_ctl_exception ;
	assign \Core_2stage.d_io_ctl_exception_cause_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_ctl_exception_cause_obs_trg_arg0 = \Core_2stage.d_io_ctl_exception_cause ;
	assign \Core_2stage.d_io_ctl_if_kill_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_ctl_if_kill_obs_trg_arg0 = \Core_2stage.d_io_ctl_if_kill ;
	assign \Core_2stage.d_io_ctl_mem_fcn_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_ctl_mem_fcn_obs_trg_arg0 = \Core_2stage.d_io_ctl_mem_fcn ;
	assign \Core_2stage.d_io_ctl_mem_typ_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_ctl_mem_typ_obs_trg_arg0 = \Core_2stage.d_io_ctl_mem_typ ;
	assign \Core_2stage.d_io_ctl_mem_val_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_ctl_mem_val_obs_trg_arg0 = \Core_2stage.d_io_ctl_mem_val ;
	assign \Core_2stage.d_io_ctl_op1_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_ctl_op1_sel_obs_trg_arg0 = \Core_2stage.d_io_ctl_op1_sel ;
	assign \Core_2stage.d_io_ctl_op2_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_ctl_op2_sel_obs_trg_arg0 = \Core_2stage.d_io_ctl_op2_sel ;
	assign \Core_2stage.d_io_ctl_pc_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_ctl_pc_sel_obs_trg_arg0 = \Core_2stage.d_io_ctl_pc_sel ;
	assign \Core_2stage.d_io_ctl_pc_sel_no_xept_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_ctl_pc_sel_no_xept_obs_trg_arg0 = \Core_2stage.d_io_ctl_pc_sel_no_xept ;
	assign \Core_2stage.d_io_ctl_rf_wen_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_ctl_rf_wen_obs_trg_arg0 = \Core_2stage.d_io_ctl_rf_wen ;
	assign \Core_2stage.d_io_ctl_stall_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_ctl_stall_obs_trg_arg0 = \Core_2stage.d_io_ctl_stall ;
	assign \Core_2stage.d_io_ctl_wb_sel_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_ctl_wb_sel_obs_trg_arg0 = \Core_2stage.d_io_ctl_wb_sel ;
	assign \Core_2stage.d_io_dat_br_eq_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_dat_br_eq_obs_trg_arg0 = \Core_2stage.d_io_dat_br_eq ;
	assign \Core_2stage.d_io_dat_br_lt_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_dat_br_lt_obs_trg_arg0 = \Core_2stage.d_io_dat_br_lt ;
	assign \Core_2stage.d_io_dat_br_ltu_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_dat_br_ltu_obs_trg_arg0 = \Core_2stage.d_io_dat_br_ltu ;
	assign \Core_2stage.d_io_dat_csr_eret_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_dat_csr_eret_obs_trg_arg0 = \Core_2stage.d_io_dat_csr_eret ;
	assign \Core_2stage.d_io_dat_csr_interrupt_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_dat_csr_interrupt_obs_trg_arg0 = \Core_2stage.d_io_dat_csr_interrupt ;
	assign \Core_2stage.d_io_dat_data_misaligned_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_dat_data_misaligned_obs_trg_arg0 = \Core_2stage.d_io_dat_data_misaligned ;
	assign \Core_2stage.d_io_dat_if_valid_resp_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_dat_if_valid_resp_obs_trg_arg0 = \Core_2stage.d_io_dat_if_valid_resp ;
	assign \Core_2stage.d_io_dat_inst_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_dat_inst_obs_trg_arg0 = \Core_2stage.d_io_dat_inst ;
	assign \Core_2stage.d_io_dat_inst_misaligned_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_dat_inst_misaligned_obs_trg_arg0 = \Core_2stage.d_io_dat_inst_misaligned ;
	assign \Core_2stage.d_io_dat_mem_store_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_dat_mem_store_obs_trg_arg0 = \Core_2stage.d_io_dat_mem_store ;
	assign \Core_2stage.d_io_dmem_req_bits_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_dmem_req_bits_addr_obs_trg_arg0 = \Core_2stage.d_io_dmem_req_bits_addr ;
	assign \Core_2stage.d_io_dmem_req_bits_data_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_dmem_req_bits_data_obs_trg_arg0 = \Core_2stage.d_io_dmem_req_bits_data ;
	assign \Core_2stage.d_io_dmem_resp_bits_data_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_dmem_resp_bits_data_obs_trg_arg0 = \Core_2stage.d_io_dmem_resp_bits_data ;
	assign \Core_2stage.d_io_hartid_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_hartid_obs_trg_arg0 = \Core_2stage.d_io_hartid ;
	assign \Core_2stage.d_io_imem_req_bits_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_imem_req_bits_addr_obs_trg_arg0 = \Core_2stage.d_io_imem_req_bits_addr ;
	assign \Core_2stage.d_io_imem_req_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_imem_req_valid_obs_trg_arg0 = \Core_2stage.d_io_imem_req_valid ;
	assign \Core_2stage.d_io_imem_resp_bits_data_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_imem_resp_bits_data_obs_trg_arg0 = \Core_2stage.d_io_imem_resp_bits_data ;
	assign \Core_2stage.d_io_imem_resp_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_imem_resp_valid_obs_trg_arg0 = \Core_2stage.d_io_imem_resp_valid ;
	assign \Core_2stage.d_io_interrupt_debug_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_interrupt_debug_obs_trg_arg0 = \Core_2stage.d_io_interrupt_debug ;
	assign \Core_2stage.d_io_interrupt_meip_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_interrupt_meip_obs_trg_arg0 = \Core_2stage.d_io_interrupt_meip ;
	assign \Core_2stage.d_io_interrupt_msip_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_interrupt_msip_obs_trg_arg0 = \Core_2stage.d_io_interrupt_msip ;
	assign \Core_2stage.d_io_interrupt_mtip_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_interrupt_mtip_obs_trg_arg0 = \Core_2stage.d_io_interrupt_mtip ;
	assign \Core_2stage.d_io_reset_vector_obs_trg_cond = 1 ;
	assign \Core_2stage.d_io_reset_vector_obs_trg_arg0 = \Core_2stage.d_io_reset_vector ;
	assign \Core_2stage.d_reset_obs_trg_cond = 1 ;
	assign \Core_2stage.d_reset_obs_trg_arg0 = \Core_2stage.d_reset ;
	assign \Core_2stage.io_dmem_req_bits_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.io_dmem_req_bits_addr_obs_trg_arg0 = \Core_2stage.io_dmem_req_bits_addr ;
	assign \Core_2stage.io_dmem_req_bits_data_obs_trg_cond = 1 ;
	assign \Core_2stage.io_dmem_req_bits_data_obs_trg_arg0 = \Core_2stage.io_dmem_req_bits_data ;
	assign \Core_2stage.io_dmem_req_bits_fcn_obs_trg_cond = 1 ;
	assign \Core_2stage.io_dmem_req_bits_fcn_obs_trg_arg0 = \Core_2stage.io_dmem_req_bits_fcn ;
	assign \Core_2stage.io_dmem_req_bits_typ_obs_trg_cond = 1 ;
	assign \Core_2stage.io_dmem_req_bits_typ_obs_trg_arg0 = \Core_2stage.io_dmem_req_bits_typ ;
	assign \Core_2stage.io_dmem_req_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.io_dmem_req_valid_obs_trg_arg0 = \Core_2stage.io_dmem_req_valid ;
	assign \Core_2stage.io_dmem_resp_bits_data_obs_trg_cond = 1 ;
	assign \Core_2stage.io_dmem_resp_bits_data_obs_trg_arg0 = \Core_2stage.io_dmem_resp_bits_data ;
	assign \Core_2stage.io_dmem_resp_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.io_dmem_resp_valid_obs_trg_arg0 = \Core_2stage.io_dmem_resp_valid ;
	assign \Core_2stage.io_hartid_obs_trg_cond = 1 ;
	assign \Core_2stage.io_hartid_obs_trg_arg0 = \Core_2stage.io_hartid ;
	assign \Core_2stage.io_imem_req_bits_addr_obs_trg_cond = 1 ;
	assign \Core_2stage.io_imem_req_bits_addr_obs_trg_arg0 = \Core_2stage.io_imem_req_bits_addr ;
	assign \Core_2stage.io_imem_req_bits_addr_state_invariant_obs_trg_cond = 1 ;
	assign \Core_2stage.io_imem_req_bits_addr_state_invariant_obs_trg_arg0 = \Core_2stage.io_imem_req_bits_addr_state_invariant ;
	assign \Core_2stage.io_imem_req_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.io_imem_req_valid_obs_trg_arg0 = \Core_2stage.io_imem_req_valid ;
	assign \Core_2stage.io_imem_resp_bits_data_obs_trg_cond = 1 ;
	assign \Core_2stage.io_imem_resp_bits_data_obs_trg_arg0 = \Core_2stage.io_imem_resp_bits_data ;
	assign \Core_2stage.io_imem_resp_bits_data_state_invariant_obs_trg_cond = 1 ;
	assign \Core_2stage.io_imem_resp_bits_data_state_invariant_obs_trg_arg0 = \Core_2stage.io_imem_resp_bits_data_state_invariant ;
	assign \Core_2stage.io_imem_resp_valid_obs_trg_cond = 1 ;
	assign \Core_2stage.io_imem_resp_valid_obs_trg_arg0 = \Core_2stage.io_imem_resp_valid ;
	assign \Core_2stage.io_interrupt_debug_obs_trg_cond = 1 ;
	assign \Core_2stage.io_interrupt_debug_obs_trg_arg0 = \Core_2stage.io_interrupt_debug ;
	assign \Core_2stage.io_interrupt_meip_obs_trg_cond = 1 ;
	assign \Core_2stage.io_interrupt_meip_obs_trg_arg0 = \Core_2stage.io_interrupt_meip ;
	assign \Core_2stage.io_interrupt_msip_obs_trg_cond = 1 ;
	assign \Core_2stage.io_interrupt_msip_obs_trg_arg0 = \Core_2stage.io_interrupt_msip ;
	assign \Core_2stage.io_interrupt_mtip_obs_trg_cond = 1 ;
	assign \Core_2stage.io_interrupt_mtip_obs_trg_arg0 = \Core_2stage.io_interrupt_mtip ;
	assign \Core_2stage.io_reset_vector_obs_trg_cond = 1 ;
	assign \Core_2stage.io_reset_vector_obs_trg_arg0 = \Core_2stage.io_reset_vector ;
	assign \Core_2stage.reset_obs_trg_cond = 1 ;
	assign \Core_2stage.reset_obs_trg_arg0 = \Core_2stage.reset ;
	assign \SodorRequestRouter_2stage_0._in_range_T_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0._in_range_T_obs_trg_arg0 = \SodorRequestRouter_2stage_0._in_range_T ;
	assign \SodorRequestRouter_2stage_0._in_range_T_1_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0._in_range_T_1_obs_trg_arg0 = \SodorRequestRouter_2stage_0._in_range_T_1 ;
	assign \SodorRequestRouter_2stage_0._in_range_T_3_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0._in_range_T_3_obs_trg_arg0 = \SodorRequestRouter_2stage_0._in_range_T_3 ;
	assign \SodorRequestRouter_2stage_0._resp_in_range_T_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0._resp_in_range_T_obs_trg_arg0 = \SodorRequestRouter_2stage_0._resp_in_range_T ;
	assign \SodorRequestRouter_2stage_0._resp_in_range_T_1_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0._resp_in_range_T_1_obs_trg_arg0 = \SodorRequestRouter_2stage_0._resp_in_range_T_1 ;
	assign \SodorRequestRouter_2stage_0._resp_in_range_T_3_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0._resp_in_range_T_3_obs_trg_arg0 = \SodorRequestRouter_2stage_0._resp_in_range_T_3 ;
	assign \SodorRequestRouter_2stage_0.in_range_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.in_range_obs_trg_arg0 = \SodorRequestRouter_2stage_0.in_range ;
	assign \SodorRequestRouter_2stage_0.io_corePort_req_bits_addr_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_corePort_req_bits_addr_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_corePort_req_bits_addr ;
	assign \SodorRequestRouter_2stage_0.io_corePort_req_bits_data_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_corePort_req_bits_data_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_corePort_req_bits_data ;
	assign \SodorRequestRouter_2stage_0.io_corePort_req_bits_fcn_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_corePort_req_bits_fcn_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_corePort_req_bits_fcn ;
	assign \SodorRequestRouter_2stage_0.io_corePort_req_bits_typ_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_corePort_req_bits_typ_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_corePort_req_bits_typ ;
	assign \SodorRequestRouter_2stage_0.io_corePort_req_valid_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_corePort_req_valid_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_corePort_req_valid ;
	assign \SodorRequestRouter_2stage_0.io_corePort_resp_bits_data_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_corePort_resp_bits_data_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_corePort_resp_bits_data ;
	assign \SodorRequestRouter_2stage_0.io_corePort_resp_valid_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_corePort_resp_valid_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_corePort_resp_valid ;
	assign \SodorRequestRouter_2stage_0.io_masterPort_req_bits_addr_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_masterPort_req_bits_addr_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_masterPort_req_bits_addr ;
	assign \SodorRequestRouter_2stage_0.io_masterPort_req_bits_data_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_masterPort_req_bits_data_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_masterPort_req_bits_data ;
	assign \SodorRequestRouter_2stage_0.io_masterPort_req_bits_fcn_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_masterPort_req_bits_fcn_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_masterPort_req_bits_fcn ;
	assign \SodorRequestRouter_2stage_0.io_masterPort_req_bits_typ_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_masterPort_req_bits_typ_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_masterPort_req_bits_typ ;
	assign \SodorRequestRouter_2stage_0.io_masterPort_req_valid_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_masterPort_req_valid_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_masterPort_req_valid ;
	assign \SodorRequestRouter_2stage_0.io_masterPort_resp_bits_data_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_masterPort_resp_bits_data_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_masterPort_resp_bits_data ;
	assign \SodorRequestRouter_2stage_0.io_masterPort_resp_valid_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_masterPort_resp_valid_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_masterPort_resp_valid ;
	assign \SodorRequestRouter_2stage_0.io_respAddress_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_respAddress_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_respAddress ;
	assign \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_addr_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_addr_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_addr ;
	assign \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_data_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_data_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_data ;
	assign \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_fcn_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_fcn_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_fcn ;
	assign \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_typ_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_typ_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_scratchPort_req_bits_typ ;
	assign \SodorRequestRouter_2stage_0.io_scratchPort_req_valid_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_scratchPort_req_valid_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_scratchPort_req_valid ;
	assign \SodorRequestRouter_2stage_0.io_scratchPort_resp_bits_data_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_scratchPort_resp_bits_data_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_scratchPort_resp_bits_data ;
	assign \SodorRequestRouter_2stage_0.io_scratchPort_resp_valid_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.io_scratchPort_resp_valid_obs_trg_arg0 = \SodorRequestRouter_2stage_0.io_scratchPort_resp_valid ;
	assign \SodorRequestRouter_2stage_0.resp_in_range_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_0.resp_in_range_obs_trg_arg0 = \SodorRequestRouter_2stage_0.resp_in_range ;
	assign \SodorRequestRouter_2stage_1._in_range_T_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1._in_range_T_obs_trg_arg0 = \SodorRequestRouter_2stage_1._in_range_T ;
	assign \SodorRequestRouter_2stage_1._in_range_T_1_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1._in_range_T_1_obs_trg_arg0 = \SodorRequestRouter_2stage_1._in_range_T_1 ;
	assign \SodorRequestRouter_2stage_1._in_range_T_3_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1._in_range_T_3_obs_trg_arg0 = \SodorRequestRouter_2stage_1._in_range_T_3 ;
	assign \SodorRequestRouter_2stage_1._resp_in_range_T_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1._resp_in_range_T_obs_trg_arg0 = \SodorRequestRouter_2stage_1._resp_in_range_T ;
	assign \SodorRequestRouter_2stage_1._resp_in_range_T_1_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1._resp_in_range_T_1_obs_trg_arg0 = \SodorRequestRouter_2stage_1._resp_in_range_T_1 ;
	assign \SodorRequestRouter_2stage_1._resp_in_range_T_3_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1._resp_in_range_T_3_obs_trg_arg0 = \SodorRequestRouter_2stage_1._resp_in_range_T_3 ;
	assign \SodorRequestRouter_2stage_1.in_range_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.in_range_obs_trg_arg0 = \SodorRequestRouter_2stage_1.in_range ;
	assign \SodorRequestRouter_2stage_1.io_corePort_req_bits_addr_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_corePort_req_bits_addr_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_corePort_req_bits_addr ;
	assign \SodorRequestRouter_2stage_1.io_corePort_req_bits_data_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_corePort_req_bits_data_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_corePort_req_bits_data ;
	assign \SodorRequestRouter_2stage_1.io_corePort_req_bits_fcn_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_corePort_req_bits_fcn_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_corePort_req_bits_fcn ;
	assign \SodorRequestRouter_2stage_1.io_corePort_req_bits_typ_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_corePort_req_bits_typ_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_corePort_req_bits_typ ;
	assign \SodorRequestRouter_2stage_1.io_corePort_req_valid_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_corePort_req_valid_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_corePort_req_valid ;
	assign \SodorRequestRouter_2stage_1.io_corePort_resp_bits_data_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_corePort_resp_bits_data_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_corePort_resp_bits_data ;
	assign \SodorRequestRouter_2stage_1.io_corePort_resp_valid_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_corePort_resp_valid_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_corePort_resp_valid ;
	assign \SodorRequestRouter_2stage_1.io_masterPort_req_bits_addr_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_masterPort_req_bits_addr_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_masterPort_req_bits_addr ;
	assign \SodorRequestRouter_2stage_1.io_masterPort_req_bits_data_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_masterPort_req_bits_data_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_masterPort_req_bits_data ;
	assign \SodorRequestRouter_2stage_1.io_masterPort_req_bits_fcn_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_masterPort_req_bits_fcn_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_masterPort_req_bits_fcn ;
	assign \SodorRequestRouter_2stage_1.io_masterPort_req_bits_typ_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_masterPort_req_bits_typ_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_masterPort_req_bits_typ ;
	assign \SodorRequestRouter_2stage_1.io_masterPort_req_valid_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_masterPort_req_valid_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_masterPort_req_valid ;
	assign \SodorRequestRouter_2stage_1.io_masterPort_resp_bits_data_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_masterPort_resp_bits_data_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_masterPort_resp_bits_data ;
	assign \SodorRequestRouter_2stage_1.io_masterPort_resp_valid_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_masterPort_resp_valid_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_masterPort_resp_valid ;
	assign \SodorRequestRouter_2stage_1.io_respAddress_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_respAddress_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_respAddress ;
	assign \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_addr_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_addr_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_addr ;
	assign \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_data_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_data_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_data ;
	assign \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_fcn_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_fcn_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_fcn ;
	assign \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_typ_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_typ_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_scratchPort_req_bits_typ ;
	assign \SodorRequestRouter_2stage_1.io_scratchPort_req_valid_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_scratchPort_req_valid_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_scratchPort_req_valid ;
	assign \SodorRequestRouter_2stage_1.io_scratchPort_resp_bits_data_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_scratchPort_resp_bits_data_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_scratchPort_resp_bits_data ;
	assign \SodorRequestRouter_2stage_1.io_scratchPort_resp_valid_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.io_scratchPort_resp_valid_obs_trg_arg0 = \SodorRequestRouter_2stage_1.io_scratchPort_resp_valid ;
	assign \SodorRequestRouter_2stage_1.resp_in_range_obs_trg_cond = 1 ;
	assign \SodorRequestRouter_2stage_1.resp_in_range_obs_trg_arg0 = \SodorRequestRouter_2stage_1.resp_in_range ;
	assign clock_obs_trg_cond = 1 ;
	assign clock_obs_trg_arg0 = clock ;
	assign core_clock_obs_trg_cond = 1 ;
	assign core_clock_obs_trg_arg0 = core_clock ;
	assign core_io_dmem_req_bits_addr_obs_trg_cond = 1 ;
	assign core_io_dmem_req_bits_addr_obs_trg_arg0 = core_io_dmem_req_bits_addr ;
	assign core_io_dmem_req_bits_data_obs_trg_cond = 1 ;
	assign core_io_dmem_req_bits_data_obs_trg_arg0 = core_io_dmem_req_bits_data ;
	assign core_io_dmem_req_bits_fcn_obs_trg_cond = 1 ;
	assign core_io_dmem_req_bits_fcn_obs_trg_arg0 = core_io_dmem_req_bits_fcn ;
	assign core_io_dmem_req_bits_typ_obs_trg_cond = 1 ;
	assign core_io_dmem_req_bits_typ_obs_trg_arg0 = core_io_dmem_req_bits_typ ;
	assign core_io_dmem_req_valid_obs_trg_cond = 1 ;
	assign core_io_dmem_req_valid_obs_trg_arg0 = core_io_dmem_req_valid ;
	assign core_io_dmem_resp_bits_data_obs_trg_cond = 1 ;
	assign core_io_dmem_resp_bits_data_obs_trg_arg0 = core_io_dmem_resp_bits_data ;
	assign core_io_dmem_resp_valid_obs_trg_cond = 1 ;
	assign core_io_dmem_resp_valid_obs_trg_arg0 = core_io_dmem_resp_valid ;
	assign core_io_hartid_obs_trg_cond = 1 ;
	assign core_io_hartid_obs_trg_arg0 = core_io_hartid ;
	assign core_io_imem_req_bits_addr_obs_trg_cond = 1 ;
	assign core_io_imem_req_bits_addr_obs_trg_arg0 = core_io_imem_req_bits_addr ;
	assign core_io_imem_req_valid_obs_trg_cond = 1 ;
	assign core_io_imem_req_valid_obs_trg_arg0 = core_io_imem_req_valid ;
	assign core_io_imem_resp_bits_data_obs_trg_cond = 1 ;
	assign core_io_imem_resp_bits_data_obs_trg_arg0 = core_io_imem_resp_bits_data ;
	assign core_io_imem_resp_valid_obs_trg_cond = 1 ;
	assign core_io_imem_resp_valid_obs_trg_arg0 = core_io_imem_resp_valid ;
	assign core_io_interrupt_debug_obs_trg_cond = 1 ;
	assign core_io_interrupt_debug_obs_trg_arg0 = core_io_interrupt_debug ;
	assign core_io_interrupt_meip_obs_trg_cond = 1 ;
	assign core_io_interrupt_meip_obs_trg_arg0 = core_io_interrupt_meip ;
	assign core_io_interrupt_msip_obs_trg_cond = 1 ;
	assign core_io_interrupt_msip_obs_trg_arg0 = core_io_interrupt_msip ;
	assign core_io_interrupt_mtip_obs_trg_cond = 1 ;
	assign core_io_interrupt_mtip_obs_trg_arg0 = core_io_interrupt_mtip ;
	assign core_io_reset_vector_obs_trg_cond = 1 ;
	assign core_io_reset_vector_obs_trg_arg0 = core_io_reset_vector ;
	assign core_reset_obs_trg_cond = 1 ;
	assign core_reset_obs_trg_arg0 = core_reset ;
	assign io_debug_port_req_bits_addr_obs_trg_cond = 1 ;
	assign io_debug_port_req_bits_addr_obs_trg_arg0 = io_debug_port_req_bits_addr ;
	assign io_debug_port_req_bits_data_obs_trg_cond = 1 ;
	assign io_debug_port_req_bits_data_obs_trg_arg0 = io_debug_port_req_bits_data ;
	assign io_debug_port_req_bits_fcn_obs_trg_cond = 1 ;
	assign io_debug_port_req_bits_fcn_obs_trg_arg0 = io_debug_port_req_bits_fcn ;
	assign io_debug_port_req_bits_typ_obs_trg_cond = 1 ;
	assign io_debug_port_req_bits_typ_obs_trg_arg0 = io_debug_port_req_bits_typ ;
	assign io_debug_port_req_valid_obs_trg_cond = 1 ;
	assign io_debug_port_req_valid_obs_trg_arg0 = io_debug_port_req_valid ;
	assign io_debug_port_resp_bits_data_obs_trg_cond = 1 ;
	assign io_debug_port_resp_bits_data_obs_trg_arg0 = io_debug_port_resp_bits_data ;
	assign io_debug_port_resp_valid_obs_trg_cond = 1 ;
	assign io_debug_port_resp_valid_obs_trg_arg0 = io_debug_port_resp_valid ;
	assign io_hartid_obs_trg_cond = 1 ;
	assign io_hartid_obs_trg_arg0 = io_hartid ;
	assign io_imem_req_bits_addr_state_invariant_obs_trg_cond = 1 ;
	assign io_imem_req_bits_addr_state_invariant_obs_trg_arg0 = io_imem_req_bits_addr_state_invariant ;
	assign io_imem_resp_bits_data_state_invariant_obs_trg_cond = 1 ;
	assign io_imem_resp_bits_data_state_invariant_obs_trg_arg0 = io_imem_resp_bits_data_state_invariant ;
	assign io_interrupt_debug_obs_trg_cond = 1 ;
	assign io_interrupt_debug_obs_trg_arg0 = io_interrupt_debug ;
	assign io_interrupt_meip_obs_trg_cond = 1 ;
	assign io_interrupt_meip_obs_trg_arg0 = io_interrupt_meip ;
	assign io_interrupt_msip_obs_trg_cond = 1 ;
	assign io_interrupt_msip_obs_trg_arg0 = io_interrupt_msip ;
	assign io_interrupt_mtip_obs_trg_cond = 1 ;
	assign io_interrupt_mtip_obs_trg_arg0 = io_interrupt_mtip ;
	assign io_master_port_0_req_bits_addr_obs_trg_cond = 1 ;
	assign io_master_port_0_req_bits_addr_obs_trg_arg0 = io_master_port_0_req_bits_addr ;
	assign io_master_port_0_req_bits_data_obs_trg_cond = 1 ;
	assign io_master_port_0_req_bits_data_obs_trg_arg0 = io_master_port_0_req_bits_data ;
	assign io_master_port_0_req_bits_fcn_obs_trg_cond = 1 ;
	assign io_master_port_0_req_bits_fcn_obs_trg_arg0 = io_master_port_0_req_bits_fcn ;
	assign io_master_port_0_req_bits_typ_obs_trg_cond = 1 ;
	assign io_master_port_0_req_bits_typ_obs_trg_arg0 = io_master_port_0_req_bits_typ ;
	assign io_master_port_0_req_valid_obs_trg_cond = 1 ;
	assign io_master_port_0_req_valid_obs_trg_arg0 = io_master_port_0_req_valid ;
	assign io_master_port_0_resp_bits_data_obs_trg_cond = 1 ;
	assign io_master_port_0_resp_bits_data_obs_trg_arg0 = io_master_port_0_resp_bits_data ;
	assign io_master_port_0_resp_valid_obs_trg_cond = 1 ;
	assign io_master_port_0_resp_valid_obs_trg_arg0 = io_master_port_0_resp_valid ;
	assign io_master_port_1_req_bits_addr_obs_trg_cond = 1 ;
	assign io_master_port_1_req_bits_addr_obs_trg_arg0 = io_master_port_1_req_bits_addr ;
	assign io_master_port_1_req_bits_data_obs_trg_cond = 1 ;
	assign io_master_port_1_req_bits_data_obs_trg_arg0 = io_master_port_1_req_bits_data ;
	assign io_master_port_1_req_bits_fcn_obs_trg_cond = 1 ;
	assign io_master_port_1_req_bits_fcn_obs_trg_arg0 = io_master_port_1_req_bits_fcn ;
	assign io_master_port_1_req_bits_typ_obs_trg_cond = 1 ;
	assign io_master_port_1_req_bits_typ_obs_trg_arg0 = io_master_port_1_req_bits_typ ;
	assign io_master_port_1_req_valid_obs_trg_cond = 1 ;
	assign io_master_port_1_req_valid_obs_trg_arg0 = io_master_port_1_req_valid ;
	assign io_master_port_1_resp_bits_data_obs_trg_cond = 1 ;
	assign io_master_port_1_resp_bits_data_obs_trg_arg0 = io_master_port_1_resp_bits_data ;
	assign io_master_port_1_resp_valid_obs_trg_cond = 1 ;
	assign io_master_port_1_resp_valid_obs_trg_arg0 = io_master_port_1_resp_valid ;
	assign io_reset_vector_obs_trg_cond = 1 ;
	assign io_reset_vector_obs_trg_arg0 = io_reset_vector ;
	assign memory_clock_obs_trg_cond = 1 ;
	assign memory_clock_obs_trg_arg0 = memory_clock ;
	assign memory_io_core_ports_0_req_bits_addr_obs_trg_cond = 1 ;
	assign memory_io_core_ports_0_req_bits_addr_obs_trg_arg0 = memory_io_core_ports_0_req_bits_addr ;
	assign memory_io_core_ports_0_req_bits_data_obs_trg_cond = 1 ;
	assign memory_io_core_ports_0_req_bits_data_obs_trg_arg0 = memory_io_core_ports_0_req_bits_data ;
	assign memory_io_core_ports_0_req_bits_fcn_obs_trg_cond = 1 ;
	assign memory_io_core_ports_0_req_bits_fcn_obs_trg_arg0 = memory_io_core_ports_0_req_bits_fcn ;
	assign memory_io_core_ports_0_req_bits_typ_obs_trg_cond = 1 ;
	assign memory_io_core_ports_0_req_bits_typ_obs_trg_arg0 = memory_io_core_ports_0_req_bits_typ ;
	assign memory_io_core_ports_0_req_valid_obs_trg_cond = 1 ;
	assign memory_io_core_ports_0_req_valid_obs_trg_arg0 = memory_io_core_ports_0_req_valid ;
	assign memory_io_core_ports_0_resp_bits_data_obs_trg_cond = 1 ;
	assign memory_io_core_ports_0_resp_bits_data_obs_trg_arg0 = memory_io_core_ports_0_resp_bits_data ;
	assign memory_io_core_ports_0_resp_valid_obs_trg_cond = 1 ;
	assign memory_io_core_ports_0_resp_valid_obs_trg_arg0 = memory_io_core_ports_0_resp_valid ;
	assign memory_io_core_ports_1_req_bits_addr_obs_trg_cond = 1 ;
	assign memory_io_core_ports_1_req_bits_addr_obs_trg_arg0 = memory_io_core_ports_1_req_bits_addr ;
	assign memory_io_core_ports_1_req_bits_typ_obs_trg_cond = 1 ;
	assign memory_io_core_ports_1_req_bits_typ_obs_trg_arg0 = memory_io_core_ports_1_req_bits_typ ;
	assign memory_io_core_ports_1_req_valid_obs_trg_cond = 1 ;
	assign memory_io_core_ports_1_req_valid_obs_trg_arg0 = memory_io_core_ports_1_req_valid ;
	assign memory_io_core_ports_1_resp_bits_data_obs_trg_cond = 1 ;
	assign memory_io_core_ports_1_resp_bits_data_obs_trg_arg0 = memory_io_core_ports_1_resp_bits_data ;
	assign memory_io_core_ports_1_resp_valid_obs_trg_cond = 1 ;
	assign memory_io_core_ports_1_resp_valid_obs_trg_arg0 = memory_io_core_ports_1_resp_valid ;
	assign memory_io_debug_port_req_bits_addr_obs_trg_cond = 1 ;
	assign memory_io_debug_port_req_bits_addr_obs_trg_arg0 = memory_io_debug_port_req_bits_addr ;
	assign memory_io_debug_port_req_bits_data_obs_trg_cond = 1 ;
	assign memory_io_debug_port_req_bits_data_obs_trg_arg0 = memory_io_debug_port_req_bits_data ;
	assign memory_io_debug_port_req_bits_fcn_obs_trg_cond = 1 ;
	assign memory_io_debug_port_req_bits_fcn_obs_trg_arg0 = memory_io_debug_port_req_bits_fcn ;
	assign memory_io_debug_port_req_bits_typ_obs_trg_cond = 1 ;
	assign memory_io_debug_port_req_bits_typ_obs_trg_arg0 = memory_io_debug_port_req_bits_typ ;
	assign memory_io_debug_port_req_valid_obs_trg_cond = 1 ;
	assign memory_io_debug_port_req_valid_obs_trg_arg0 = memory_io_debug_port_req_valid ;
	assign memory_io_debug_port_resp_bits_data_obs_trg_cond = 1 ;
	assign memory_io_debug_port_resp_bits_data_obs_trg_arg0 = memory_io_debug_port_resp_bits_data ;
	assign memory_io_debug_port_resp_valid_obs_trg_cond = 1 ;
	assign memory_io_debug_port_resp_valid_obs_trg_arg0 = memory_io_debug_port_resp_valid ;
	assign reset_obs_trg_cond = 1 ;
	assign reset_obs_trg_arg0 = reset ;
	assign router_1_io_corePort_req_bits_addr_obs_trg_cond = 1 ;
	assign router_1_io_corePort_req_bits_addr_obs_trg_arg0 = router_1_io_corePort_req_bits_addr ;
	assign router_1_io_corePort_req_bits_data_obs_trg_cond = 1 ;
	assign router_1_io_corePort_req_bits_data_obs_trg_arg0 = router_1_io_corePort_req_bits_data ;
	assign router_1_io_corePort_req_bits_fcn_obs_trg_cond = 1 ;
	assign router_1_io_corePort_req_bits_fcn_obs_trg_arg0 = router_1_io_corePort_req_bits_fcn ;
	assign router_1_io_corePort_req_bits_typ_obs_trg_cond = 1 ;
	assign router_1_io_corePort_req_bits_typ_obs_trg_arg0 = router_1_io_corePort_req_bits_typ ;
	assign router_1_io_corePort_req_valid_obs_trg_cond = 1 ;
	assign router_1_io_corePort_req_valid_obs_trg_arg0 = router_1_io_corePort_req_valid ;
	assign router_1_io_corePort_resp_bits_data_obs_trg_cond = 1 ;
	assign router_1_io_corePort_resp_bits_data_obs_trg_arg0 = router_1_io_corePort_resp_bits_data ;
	assign router_1_io_corePort_resp_valid_obs_trg_cond = 1 ;
	assign router_1_io_corePort_resp_valid_obs_trg_arg0 = router_1_io_corePort_resp_valid ;
	assign router_1_io_masterPort_req_bits_addr_obs_trg_cond = 1 ;
	assign router_1_io_masterPort_req_bits_addr_obs_trg_arg0 = router_1_io_masterPort_req_bits_addr ;
	assign router_1_io_masterPort_req_bits_data_obs_trg_cond = 1 ;
	assign router_1_io_masterPort_req_bits_data_obs_trg_arg0 = router_1_io_masterPort_req_bits_data ;
	assign router_1_io_masterPort_req_bits_fcn_obs_trg_cond = 1 ;
	assign router_1_io_masterPort_req_bits_fcn_obs_trg_arg0 = router_1_io_masterPort_req_bits_fcn ;
	assign router_1_io_masterPort_req_bits_typ_obs_trg_cond = 1 ;
	assign router_1_io_masterPort_req_bits_typ_obs_trg_arg0 = router_1_io_masterPort_req_bits_typ ;
	assign router_1_io_masterPort_req_valid_obs_trg_cond = 1 ;
	assign router_1_io_masterPort_req_valid_obs_trg_arg0 = router_1_io_masterPort_req_valid ;
	assign router_1_io_masterPort_resp_bits_data_obs_trg_cond = 1 ;
	assign router_1_io_masterPort_resp_bits_data_obs_trg_arg0 = router_1_io_masterPort_resp_bits_data ;
	assign router_1_io_masterPort_resp_valid_obs_trg_cond = 1 ;
	assign router_1_io_masterPort_resp_valid_obs_trg_arg0 = router_1_io_masterPort_resp_valid ;
	assign router_1_io_respAddress_obs_trg_cond = 1 ;
	assign router_1_io_respAddress_obs_trg_arg0 = router_1_io_respAddress ;
	assign router_1_io_scratchPort_req_bits_addr_obs_trg_cond = 1 ;
	assign router_1_io_scratchPort_req_bits_addr_obs_trg_arg0 = router_1_io_scratchPort_req_bits_addr ;
	assign router_1_io_scratchPort_req_bits_data_obs_trg_cond = 1 ;
	assign router_1_io_scratchPort_req_bits_data_obs_trg_arg0 = router_1_io_scratchPort_req_bits_data ;
	assign router_1_io_scratchPort_req_bits_fcn_obs_trg_cond = 1 ;
	assign router_1_io_scratchPort_req_bits_fcn_obs_trg_arg0 = router_1_io_scratchPort_req_bits_fcn ;
	assign router_1_io_scratchPort_req_bits_typ_obs_trg_cond = 1 ;
	assign router_1_io_scratchPort_req_bits_typ_obs_trg_arg0 = router_1_io_scratchPort_req_bits_typ ;
	assign router_1_io_scratchPort_req_valid_obs_trg_cond = 1 ;
	assign router_1_io_scratchPort_req_valid_obs_trg_arg0 = router_1_io_scratchPort_req_valid ;
	assign router_1_io_scratchPort_resp_bits_data_obs_trg_cond = 1 ;
	assign router_1_io_scratchPort_resp_bits_data_obs_trg_arg0 = router_1_io_scratchPort_resp_bits_data ;
	assign router_1_io_scratchPort_resp_valid_obs_trg_cond = 1 ;
	assign router_1_io_scratchPort_resp_valid_obs_trg_arg0 = router_1_io_scratchPort_resp_valid ;
	assign router_io_corePort_req_bits_addr_obs_trg_cond = 1 ;
	assign router_io_corePort_req_bits_addr_obs_trg_arg0 = router_io_corePort_req_bits_addr ;
	assign router_io_corePort_req_bits_data_obs_trg_cond = 1 ;
	assign router_io_corePort_req_bits_data_obs_trg_arg0 = router_io_corePort_req_bits_data ;
	assign router_io_corePort_req_bits_fcn_obs_trg_cond = 1 ;
	assign router_io_corePort_req_bits_fcn_obs_trg_arg0 = router_io_corePort_req_bits_fcn ;
	assign router_io_corePort_req_bits_typ_obs_trg_cond = 1 ;
	assign router_io_corePort_req_bits_typ_obs_trg_arg0 = router_io_corePort_req_bits_typ ;
	assign router_io_corePort_req_valid_obs_trg_cond = 1 ;
	assign router_io_corePort_req_valid_obs_trg_arg0 = router_io_corePort_req_valid ;
	assign router_io_corePort_resp_bits_data_obs_trg_cond = 1 ;
	assign router_io_corePort_resp_bits_data_obs_trg_arg0 = router_io_corePort_resp_bits_data ;
	assign router_io_corePort_resp_valid_obs_trg_cond = 1 ;
	assign router_io_corePort_resp_valid_obs_trg_arg0 = router_io_corePort_resp_valid ;
	assign router_io_masterPort_req_bits_addr_obs_trg_cond = 1 ;
	assign router_io_masterPort_req_bits_addr_obs_trg_arg0 = router_io_masterPort_req_bits_addr ;
	assign router_io_masterPort_req_bits_data_obs_trg_cond = 1 ;
	assign router_io_masterPort_req_bits_data_obs_trg_arg0 = router_io_masterPort_req_bits_data ;
	assign router_io_masterPort_req_bits_fcn_obs_trg_cond = 1 ;
	assign router_io_masterPort_req_bits_fcn_obs_trg_arg0 = router_io_masterPort_req_bits_fcn ;
	assign router_io_masterPort_req_bits_typ_obs_trg_cond = 1 ;
	assign router_io_masterPort_req_bits_typ_obs_trg_arg0 = router_io_masterPort_req_bits_typ ;
	assign router_io_masterPort_req_valid_obs_trg_cond = 1 ;
	assign router_io_masterPort_req_valid_obs_trg_arg0 = router_io_masterPort_req_valid ;
	assign router_io_masterPort_resp_bits_data_obs_trg_cond = 1 ;
	assign router_io_masterPort_resp_bits_data_obs_trg_arg0 = router_io_masterPort_resp_bits_data ;
	assign router_io_masterPort_resp_valid_obs_trg_cond = 1 ;
	assign router_io_masterPort_resp_valid_obs_trg_arg0 = router_io_masterPort_resp_valid ;
	assign router_io_respAddress_obs_trg_cond = 1 ;
	assign router_io_respAddress_obs_trg_arg0 = router_io_respAddress ;
	assign router_io_scratchPort_req_bits_addr_obs_trg_cond = 1 ;
	assign router_io_scratchPort_req_bits_addr_obs_trg_arg0 = router_io_scratchPort_req_bits_addr ;
	assign router_io_scratchPort_req_bits_data_obs_trg_cond = 1 ;
	assign router_io_scratchPort_req_bits_data_obs_trg_arg0 = router_io_scratchPort_req_bits_data ;
	assign router_io_scratchPort_req_bits_fcn_obs_trg_cond = 1 ;
	assign router_io_scratchPort_req_bits_fcn_obs_trg_arg0 = router_io_scratchPort_req_bits_fcn ;
	assign router_io_scratchPort_req_bits_typ_obs_trg_cond = 1 ;
	assign router_io_scratchPort_req_bits_typ_obs_trg_arg0 = router_io_scratchPort_req_bits_typ ;
	assign router_io_scratchPort_req_valid_obs_trg_cond = 1 ;
	assign router_io_scratchPort_req_valid_obs_trg_arg0 = router_io_scratchPort_req_valid ;
	assign router_io_scratchPort_resp_bits_data_obs_trg_cond = 1 ;
	assign router_io_scratchPort_resp_bits_data_obs_trg_arg0 = router_io_scratchPort_resp_bits_data ;
	assign router_io_scratchPort_resp_valid_obs_trg_cond = 1 ;
	assign router_io_scratchPort_resp_valid_obs_trg_arg0 = router_io_scratchPort_resp_valid ;
endmodule