module prod
(
  input clk, 
);

// Todo: defined all the wires for two copies of the circuits


//**Wire declarations**//
//**Init register**//
//**Stuttering Signal**//
//**Self-composed modules**//
//**Initial state**//
//**State invariants**//
//**Verification conditions**//

endmodule