module SodorInternalTile_2stage_state_trg ( input [31:0] \Core_2stage.DatPath_2stage.if_reg_pc , input [8191:0] mem_2_1_flat_trg , input [1023:0] regfile_flat_trg , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mpie , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_singleStepped , input [8191:0] mem_2_0_flat_trg , input [5:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.small_1 , input \Core_2stage.DatPath_2stage.reg_interrupt_handled , input [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.large_1 , input [8191:0] mem_1_1_flat_trg , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dpc , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mie , input [8191:0] mem_3_0_flat_trg , input [31:0] \Core_2stage.DatPath_2stage.if_inst_buffer , input \Core_2stage.DatPath_2stage.io_ctl_if_kill_r , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mepc , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mscratch , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mie , input [5:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.small_ , input [8191:0] mem_0_0_flat_trg , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_step , input \Core_2stage.DatPath_2stage.if_inst_buffer_valid , input [31:0] \Core_2stage.DatPath_2stage.exe_reg_pc_plus4 , input [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcountinhibit , input [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.large_ , input [8191:0] mem_0_1_flat_trg , input [31:0] \Core_2stage.DatPath_2stage.pc_x , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_debug , input [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_cause , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_wfi , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dscratch , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease_r , input [31:0] \Core_2stage.DatPath_2stage.exe_reg_pc , input \Core_2stage.DatPath_2stage.exe_reg_valid , input [8191:0] mem_3_1_flat_trg , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtval , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtvec , input [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcause , input [8191:0] mem_1_0_flat_trg , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_ebreakm , input \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_spp , input [31:0] \Core_2stage.DatPath_2stage.exe_reg_inst , output [5:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.small_1_state_trg , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtval_state_trg , output [31:0] \Core_2stage.DatPath_2stage.exe_reg_pc_state_trg , output [31:0] \Core_2stage.DatPath_2stage.exe_reg_pc_plus4_state_trg , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dpc_state_trg , output [8191:0] mem_1_1_state_trg , output [1023:0] regfile_state_trg , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcause_state_trg , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dscratch_state_trg , output \Core_2stage.DatPath_2stage.exe_reg_valid_state_trg , output [31:0] \Core_2stage.DatPath_2stage.if_reg_pc_state_trg , output [8191:0] mem_0_1_state_trg , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_ebreakm_state_trg , output [8191:0] mem_3_1_state_trg , output [8191:0] mem_3_0_state_trg , output [31:0] \Core_2stage.DatPath_2stage.if_inst_buffer_state_trg , output [5:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.small__state_trg , output \Core_2stage.DatPath_2stage.reg_interrupt_handled_state_trg , output \Core_2stage.DatPath_2stage.io_ctl_if_kill_r_state_trg , output [8191:0] mem_1_0_state_trg , output [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcountinhibit_state_trg , output \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease_r_state_trg , output [8191:0] mem_2_1_state_trg , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mscratch_state_trg , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_step_state_trg , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mie_state_trg , output [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.large_1_state_trg , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_singleStepped_state_trg , output [2:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_cause_state_trg , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_spp_state_trg , output [57:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.large__state_trg , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtvec_state_trg , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_debug_state_trg , output [31:0] \Core_2stage.DatPath_2stage.pc_x_state_trg , output \Core_2stage.DatPath_2stage.if_inst_buffer_valid_state_trg , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_wfi_state_trg , output \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mpie_state_trg , output [8191:0] mem_2_0_state_trg , output [31:0] \Core_2stage.DatPath_2stage.exe_reg_inst_state_trg , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mie_state_trg , output [31:0] \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mepc_state_trg , output [8191:0] mem_0_0_state_trg );
	assign mem_0_1_state_trg = mem_0_1_flat_trg ;
	assign mem_1_1_state_trg = mem_1_1_flat_trg ;
	assign mem_2_1_state_trg = mem_2_1_flat_trg ;
	assign mem_3_1_state_trg = mem_3_1_flat_trg ;
	assign mem_0_0_state_trg = mem_0_0_flat_trg ;
	assign mem_1_0_state_trg = mem_1_0_flat_trg ;
	assign mem_2_0_state_trg = mem_2_0_flat_trg ;
	assign mem_3_0_state_trg = mem_3_0_flat_trg ;
	assign regfile_state_trg = regfile_flat_trg ;
	assign \Core_2stage.DatPath_2stage.if_inst_buffer_state_trg = \Core_2stage.DatPath_2stage.if_inst_buffer ;
	assign \Core_2stage.DatPath_2stage.if_reg_pc_state_trg = \Core_2stage.DatPath_2stage.if_reg_pc ;
	assign \Core_2stage.DatPath_2stage.exe_reg_pc_state_trg = \Core_2stage.DatPath_2stage.exe_reg_pc ;
	assign \Core_2stage.DatPath_2stage.exe_reg_pc_plus4_state_trg = \Core_2stage.DatPath_2stage.exe_reg_pc_plus4 ;
	assign \Core_2stage.DatPath_2stage.exe_reg_inst_state_trg = \Core_2stage.DatPath_2stage.exe_reg_inst ;
	assign \Core_2stage.DatPath_2stage.exe_reg_valid_state_trg = \Core_2stage.DatPath_2stage.exe_reg_valid ;
	assign \Core_2stage.DatPath_2stage.if_inst_buffer_valid_state_trg = \Core_2stage.DatPath_2stage.if_inst_buffer_valid ;
	assign \Core_2stage.DatPath_2stage.reg_interrupt_handled_state_trg = \Core_2stage.DatPath_2stage.reg_interrupt_handled ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_wfi_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_wfi ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.small_1_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.small_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.large_1_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.large_1 ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_spp_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_spp ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mpie_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mpie ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mie_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mstatus_mie ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_ebreakm_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_ebreakm ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_cause_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_cause ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_step_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dcsr_step ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_debug_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_debug ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dpc_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dpc ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dscratch_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_dscratch ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_singleStepped_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_singleStepped ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mie_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mie ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mepc_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mepc ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcause_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcause ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtval_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtval ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mscratch_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mscratch ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtvec_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mtvec ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcountinhibit_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.reg_mcountinhibit ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.small__state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.small_ ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.large__state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.large_ ;
	assign \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease_r_state_trg = \Core_2stage.DatPath_2stage.CSRFile_2stage.io_status_cease_r ;
	assign \Core_2stage.DatPath_2stage.io_ctl_if_kill_r_state_trg = \Core_2stage.DatPath_2stage.io_ctl_if_kill_r ;
	assign \Core_2stage.DatPath_2stage.pc_x_state_trg = \Core_2stage.DatPath_2stage.pc_x ;
endmodule