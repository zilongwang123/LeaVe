module ibex_csr (
	clk_i,
	rst_ni,
	wr_data_i,
	wr_en_i,
	rd_data_o,
	rd_error_o
);
	parameter [31:0] Width = 32;
	parameter [0:0] ShadowCopy = 1'b0;
	parameter [Width - 1:0] ResetValue = 1'sb0;
	input wire clk_i;
	input wire rst_ni;
	input wire [Width - 1:0] wr_data_i;
	input wire wr_en_i;
	output wire [Width - 1:0] rd_data_o;
	output wire rd_error_o;
	reg [Width - 1:0] rdata_q;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			rdata_q <= ResetValue;
		else if (wr_en_i)
			rdata_q <= wr_data_i;
	assign rd_data_o = rdata_q;
	// generate
	// 	if (ShadowCopy) begin : gen_shadow
	// 		reg [Width - 1:0] shadow_q;
	// 		always @(posedge clk_i or negedge rst_ni)
	// 			if (!rst_ni)
	// 				shadow_q <= ~ResetValue;
	// 			else if (wr_en_i)
	// 				shadow_q <= ~wr_data_i;
	// 		assign rd_error_o = rdata_q != ~shadow_q;
	// 	end
	// 	else begin : gen_no_shadow
			assign rd_error_o = 1'b0;
	// 	end
	// endgenerate
endmodule
