module SodorInternalTile_1stage_state_src ( input [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mepc , input \Core_1stage.CtlPath_1stage.reg_mem_en , input [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mie , input [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dscratch , input [8191:0] mem_3_1_flat_src , input [1023:0] regfile_flat_src , input \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dcsr_ebreakm , input \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_singleStepped , input [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mcause , input [8191:0] mem_0_1_flat_src , input \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_wfi , input [8191:0] mem_1_0_flat_src , input [8191:0] mem_0_0_flat_src , input \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mstatus_spp , input [5:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.small_ , input [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mtval , input [2:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mcountinhibit , input \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mstatus_mpie , input [57:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.large_1 , input [8191:0] mem_1_1_flat_src , input [31:0] \Core_1stage.DatPath_1stage.if_inst_buffer , input [5:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.small_1 , input \Core_1stage.DatPath_1stage.reg_interrupt_edge , input [57:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.large_ , input [2:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dcsr_cause , input [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dpc , input [8191:0] mem_2_1_flat_src , input [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mscratch , input [31:0] \Core_1stage.DatPath_1stage.pc_reg , input [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mtvec , input \Core_1stage.DatPath_1stage.CSRFile_1stage.io_status_cease_r , input \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dcsr_step , input \Core_1stage.DatPath_1stage.reg_dmiss , input [8191:0] mem_3_0_flat_src , input \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_debug , input \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mstatus_mie , input [8191:0] mem_2_0_flat_src , output \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mstatus_mie_state_src , output \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mstatus_spp_state_src , output [8191:0] mem_0_0_state_src , output [1023:0] regfile_state_src , output [5:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.small__state_src , output [31:0] \Core_1stage.DatPath_1stage.if_inst_buffer_state_src , output \Core_1stage.DatPath_1stage.reg_interrupt_edge_state_src , output \Core_1stage.DatPath_1stage.CSRFile_1stage.io_status_cease_r_state_src , output [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mie_state_src , output [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mtval_state_src , output \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dcsr_step_state_src , output [8191:0] mem_2_0_state_src , output [2:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dcsr_cause_state_src , output \Core_1stage.DatPath_1stage.reg_dmiss_state_src , output [8191:0] mem_3_0_state_src , output [57:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.large__state_src , output [5:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.small_1_state_src , output \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dcsr_ebreakm_state_src , output \Core_1stage.CtlPath_1stage.reg_mem_en_state_src , output [8191:0] mem_1_1_state_src , output [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dpc_state_src , output \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_wfi_state_src , output \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_debug_state_src , output [57:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.large_1_state_src , output \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_singleStepped_state_src , output \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mstatus_mpie_state_src , output [8191:0] mem_2_1_state_src , output [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mepc_state_src , output [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dscratch_state_src , output [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mscratch_state_src , output [31:0] \Core_1stage.DatPath_1stage.pc_reg_state_src , output [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mcause_state_src , output [31:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mtvec_state_src , output [8191:0] mem_3_1_state_src , output [8191:0] mem_1_0_state_src , output [8191:0] mem_0_1_state_src , output [2:0] \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mcountinhibit_state_src );
	assign mem_0_1_state_src = mem_0_1_flat_src ;
	assign mem_1_1_state_src = mem_1_1_flat_src ;
	assign mem_2_1_state_src = mem_2_1_flat_src ;
	assign mem_3_1_state_src = mem_3_1_flat_src ;
	assign mem_0_0_state_src = mem_0_0_flat_src ;
	assign mem_1_0_state_src = mem_1_0_flat_src ;
	assign mem_2_0_state_src = mem_2_0_flat_src ;
	assign mem_3_0_state_src = mem_3_0_flat_src ;
	assign regfile_state_src = regfile_flat_src ;
	assign \Core_1stage.DatPath_1stage.pc_reg_state_src = \Core_1stage.DatPath_1stage.pc_reg ;
	assign \Core_1stage.DatPath_1stage.reg_dmiss_state_src = \Core_1stage.DatPath_1stage.reg_dmiss ;
	assign \Core_1stage.DatPath_1stage.if_inst_buffer_state_src = \Core_1stage.DatPath_1stage.if_inst_buffer ;
	assign \Core_1stage.DatPath_1stage.reg_interrupt_edge_state_src = \Core_1stage.DatPath_1stage.reg_interrupt_edge ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mstatus_spp_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mstatus_spp ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mstatus_mpie_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mstatus_mpie ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mstatus_mie_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mstatus_mie ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dcsr_ebreakm_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dcsr_ebreakm ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dcsr_cause_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dcsr_cause ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dcsr_step_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dcsr_step ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_debug_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_debug ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dpc_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dpc ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dscratch_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_dscratch ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_singleStepped_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_singleStepped ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mie_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mie ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mepc_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mepc ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mcause_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mcause ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mtval_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mtval ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mscratch_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mscratch ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mtvec_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mtvec ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_wfi_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_wfi ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mcountinhibit_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.reg_mcountinhibit ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.small__state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.small_ ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.large__state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.large_ ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.small_1_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.small_1 ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.large_1_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.large_1 ;
	assign \Core_1stage.DatPath_1stage.CSRFile_1stage.io_status_cease_r_state_src = \Core_1stage.DatPath_1stage.CSRFile_1stage.io_status_cease_r ;
	assign \Core_1stage.CtlPath_1stage.reg_mem_en_state_src = \Core_1stage.CtlPath_1stage.reg_mem_en ;
endmodule