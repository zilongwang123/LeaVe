module AsyncScratchPadMemory_1stage(
  input         clock,
  input         io_core_ports_0_req_valid,
  input  [31:0] io_core_ports_0_req_bits_addr,
  input  [31:0] io_core_ports_0_req_bits_data,
  input         io_core_ports_0_req_bits_fcn,
  input  [2:0]  io_core_ports_0_req_bits_typ,
  output        io_core_ports_0_resp_valid,
  output [31:0] io_core_ports_0_resp_bits_data,
  input         io_core_ports_1_req_valid,
  input  [31:0] io_core_ports_1_req_bits_addr,
  input  [2:0]  io_core_ports_1_req_bits_typ,
  output        io_core_ports_1_resp_valid,
  output [31:0] io_core_ports_1_resp_bits_data,
  input         io_debug_port_req_valid,
  input  [31:0] io_debug_port_req_bits_addr,
  input  [31:0] io_debug_port_req_bits_data,
  input         io_debug_port_req_bits_fcn,
  input  [2:0]  io_debug_port_req_bits_typ,
  output        io_debug_port_resp_valid,
  output [31:0] io_debug_port_resp_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
  reg [7:0] mem_0_0 [0:1023]; // @[memory.scala 73:31]
  reg [7:0] mem_0_1 [0:1023]; // @[memory.scala 73:31]
  wire  mem_0_io_core_ports_0_resp_bits_data_MPORT_en; // @[memory.scala 73:31]
  wire [9:0] mem_0_io_core_ports_0_resp_bits_data_MPORT_addr; // @[memory.scala 73:31]
  wire [7:0] mem_0_io_core_ports_0_resp_bits_data_MPORT_data; // @[memory.scala 73:31]
  wire  mem_0_io_core_ports_1_resp_bits_data_MPORT_en; // @[memory.scala 73:31]
  wire [9:0] mem_0_io_core_ports_1_resp_bits_data_MPORT_addr; // @[memory.scala 73:31]
  wire [7:0] mem_0_io_core_ports_1_resp_bits_data_MPORT_data; // @[memory.scala 73:31]
  wire  mem_0_io_debug_port_resp_bits_data_MPORT_en; // @[memory.scala 73:31]
  wire [9:0] mem_0_io_debug_port_resp_bits_data_MPORT_addr; // @[memory.scala 73:31]
  wire [7:0] mem_0_io_debug_port_resp_bits_data_MPORT_data; // @[memory.scala 73:31]
  wire [7:0] mem_0_MPORT_data; // @[memory.scala 73:31]
  wire [9:0] mem_0_MPORT_addr; // @[memory.scala 73:31]
  wire  mem_0_MPORT_mask; // @[memory.scala 73:31]
  wire  mem_0_MPORT_en; // @[memory.scala 73:31]
  wire [7:0] mem_0_MPORT_1_data; // @[memory.scala 73:31]
  wire [9:0] mem_0_MPORT_1_addr; // @[memory.scala 73:31]
  wire  mem_0_MPORT_1_mask; // @[memory.scala 73:31]
  wire  mem_0_MPORT_1_en; // @[memory.scala 73:31]
  reg [7:0] mem_1_0 [0:1023]; // @[memory.scala 73:31]
  reg [7:0] mem_1_1 [0:1023]; // @[memory.scala 73:31]
  wire  mem_1_io_core_ports_0_resp_bits_data_MPORT_en; // @[memory.scala 73:31]
  wire [9:0] mem_1_io_core_ports_0_resp_bits_data_MPORT_addr; // @[memory.scala 73:31]
  wire [7:0] mem_1_io_core_ports_0_resp_bits_data_MPORT_data; // @[memory.scala 73:31]
  wire  mem_1_io_core_ports_1_resp_bits_data_MPORT_en; // @[memory.scala 73:31]
  wire [9:0] mem_1_io_core_ports_1_resp_bits_data_MPORT_addr; // @[memory.scala 73:31]
  wire [7:0] mem_1_io_core_ports_1_resp_bits_data_MPORT_data; // @[memory.scala 73:31]
  wire  mem_1_io_debug_port_resp_bits_data_MPORT_en; // @[memory.scala 73:31]
  wire [9:0] mem_1_io_debug_port_resp_bits_data_MPORT_addr; // @[memory.scala 73:31]
  wire [7:0] mem_1_io_debug_port_resp_bits_data_MPORT_data; // @[memory.scala 73:31]
  wire [7:0] mem_1_MPORT_data; // @[memory.scala 73:31]
  wire [9:0] mem_1_MPORT_addr; // @[memory.scala 73:31]
  wire  mem_1_MPORT_mask; // @[memory.scala 73:31]
  wire  mem_1_MPORT_en; // @[memory.scala 73:31]
  wire [7:0] mem_1_MPORT_1_data; // @[memory.scala 73:31]
  wire [9:0] mem_1_MPORT_1_addr; // @[memory.scala 73:31]
  wire  mem_1_MPORT_1_mask; // @[memory.scala 73:31]
  wire  mem_1_MPORT_1_en; // @[memory.scala 73:31]
  reg [7:0] mem_2_0 [0:1023]; // @[memory.scala 73:31]
  reg [7:0] mem_2_1 [0:1023]; // @[memory.scala 73:31]
  wire  mem_2_io_core_ports_0_resp_bits_data_MPORT_en; // @[memory.scala 73:31]
  wire [9:0] mem_2_io_core_ports_0_resp_bits_data_MPORT_addr; // @[memory.scala 73:31]
  wire [7:0] mem_2_io_core_ports_0_resp_bits_data_MPORT_data; // @[memory.scala 73:31]
  wire  mem_2_io_core_ports_1_resp_bits_data_MPORT_en; // @[memory.scala 73:31]
  wire [9:0] mem_2_io_core_ports_1_resp_bits_data_MPORT_addr; // @[memory.scala 73:31]
  wire [7:0] mem_2_io_core_ports_1_resp_bits_data_MPORT_data; // @[memory.scala 73:31]
  wire  mem_2_io_debug_port_resp_bits_data_MPORT_en; // @[memory.scala 73:31]
  wire [9:0] mem_2_io_debug_port_resp_bits_data_MPORT_addr; // @[memory.scala 73:31]
  wire [7:0] mem_2_io_debug_port_resp_bits_data_MPORT_data; // @[memory.scala 73:31]
  wire [7:0] mem_2_MPORT_data; // @[memory.scala 73:31]
  wire [9:0] mem_2_MPORT_addr; // @[memory.scala 73:31]
  wire  mem_2_MPORT_mask; // @[memory.scala 73:31]
  wire  mem_2_MPORT_en; // @[memory.scala 73:31]
  wire [7:0] mem_2_MPORT_1_data; // @[memory.scala 73:31]
  wire [9:0] mem_2_MPORT_1_addr; // @[memory.scala 73:31]
  wire  mem_2_MPORT_1_mask; // @[memory.scala 73:31]
  wire  mem_2_MPORT_1_en; // @[memory.scala 73:31]
  reg [7:0] mem_3_0 [0:1023]; // @[memory.scala 73:31]
  reg [7:0] mem_3_1 [0:1023]; // @[memory.scala 73:31]
  wire  mem_3_io_core_ports_0_resp_bits_data_MPORT_en; // @[memory.scala 73:31]
  wire [9:0] mem_3_io_core_ports_0_resp_bits_data_MPORT_addr; // @[memory.scala 73:31]
  wire [7:0] mem_3_io_core_ports_0_resp_bits_data_MPORT_data; // @[memory.scala 73:31]
  wire  mem_3_io_core_ports_1_resp_bits_data_MPORT_en; // @[memory.scala 73:31]
  wire [9:0] mem_3_io_core_ports_1_resp_bits_data_MPORT_addr; // @[memory.scala 73:31]
  wire [7:0] mem_3_io_core_ports_1_resp_bits_data_MPORT_data; // @[memory.scala 73:31]
  wire  mem_3_io_debug_port_resp_bits_data_MPORT_en; // @[memory.scala 73:31]
  wire [9:0] mem_3_io_debug_port_resp_bits_data_MPORT_addr; // @[memory.scala 73:31]
  wire [7:0] mem_3_io_debug_port_resp_bits_data_MPORT_data; // @[memory.scala 73:31]
  wire [7:0] mem_3_MPORT_data; // @[memory.scala 73:31]
  wire [9:0] mem_3_MPORT_addr; // @[memory.scala 73:31]
  wire  mem_3_MPORT_mask; // @[memory.scala 73:31]
  wire  mem_3_MPORT_en; // @[memory.scala 73:31]
  wire [7:0] mem_3_MPORT_1_data; // @[memory.scala 73:31]
  wire [9:0] mem_3_MPORT_1_addr; // @[memory.scala 73:31]
  wire  mem_3_MPORT_1_mask; // @[memory.scala 73:31]
  wire  mem_3_MPORT_1_en; // @[memory.scala 73:31]
  wire [20:0] io_core_ports_0_resp_bits_data_module_io_addr; // @[memory.scala 120:26]
  wire [1:0] io_core_ports_0_resp_bits_data_module_io_size; // @[memory.scala 120:26]
  wire  io_core_ports_0_resp_bits_data_module_io_signed; // @[memory.scala 120:26]
  wire [31:0] io_core_ports_0_resp_bits_data_module_io_data; // @[memory.scala 120:26]
  wire [9:0] io_core_ports_0_resp_bits_data_module_io_mem_addr; // @[memory.scala 120:26]
  wire [7:0] io_core_ports_0_resp_bits_data_module_io_mem_data_0; // @[memory.scala 120:26]
  wire [7:0] io_core_ports_0_resp_bits_data_module_io_mem_data_1; // @[memory.scala 120:26]
  wire [7:0] io_core_ports_0_resp_bits_data_module_io_mem_data_2; // @[memory.scala 120:26]
  wire [7:0] io_core_ports_0_resp_bits_data_module_io_mem_data_3; // @[memory.scala 120:26]
  wire [20:0] module__io_addr; // @[memory.scala 156:26]
  wire [31:0] module__io_data; // @[memory.scala 156:26]
  wire [1:0] module__io_size; // @[memory.scala 156:26]
  wire  module__io_en; // @[memory.scala 156:26]
  wire [9:0] module__io_mem_addr; // @[memory.scala 156:26]
  wire [7:0] module__io_mem_data_0; // @[memory.scala 156:26]
  wire [7:0] module__io_mem_data_1; // @[memory.scala 156:26]
  wire [7:0] module__io_mem_data_2; // @[memory.scala 156:26]
  wire [7:0] module__io_mem_data_3; // @[memory.scala 156:26]
  wire  module__io_mem_masks_0; // @[memory.scala 156:26]
  wire  module__io_mem_masks_1; // @[memory.scala 156:26]
  wire  module__io_mem_masks_2; // @[memory.scala 156:26]
  wire  module__io_mem_masks_3; // @[memory.scala 156:26]
  wire [20:0] io_core_ports_1_resp_bits_data_module_io_addr; // @[memory.scala 120:26]
  wire [1:0] io_core_ports_1_resp_bits_data_module_io_size; // @[memory.scala 120:26]
  wire  io_core_ports_1_resp_bits_data_module_io_signed; // @[memory.scala 120:26]
  wire [31:0] io_core_ports_1_resp_bits_data_module_io_data; // @[memory.scala 120:26]
  wire [9:0] io_core_ports_1_resp_bits_data_module_io_mem_addr; // @[memory.scala 120:26]
  wire [7:0] io_core_ports_1_resp_bits_data_module_io_mem_data_0; // @[memory.scala 120:26]
  wire [7:0] io_core_ports_1_resp_bits_data_module_io_mem_data_1; // @[memory.scala 120:26]
  wire [7:0] io_core_ports_1_resp_bits_data_module_io_mem_data_2; // @[memory.scala 120:26]
  wire [7:0] io_core_ports_1_resp_bits_data_module_io_mem_data_3; // @[memory.scala 120:26]
  wire [20:0] io_debug_port_resp_bits_data_module_io_addr; // @[memory.scala 120:26]
  wire [1:0] io_debug_port_resp_bits_data_module_io_size; // @[memory.scala 120:26]
  wire  io_debug_port_resp_bits_data_module_io_signed; // @[memory.scala 120:26]
  wire [31:0] io_debug_port_resp_bits_data_module_io_data; // @[memory.scala 120:26]
  wire [9:0] io_debug_port_resp_bits_data_module_io_mem_addr; // @[memory.scala 120:26]
  wire [7:0] io_debug_port_resp_bits_data_module_io_mem_data_0; // @[memory.scala 120:26]
  wire [7:0] io_debug_port_resp_bits_data_module_io_mem_data_1; // @[memory.scala 120:26]
  wire [7:0] io_debug_port_resp_bits_data_module_io_mem_data_2; // @[memory.scala 120:26]
  wire [7:0] io_debug_port_resp_bits_data_module_io_mem_data_3; // @[memory.scala 120:26]
  wire [20:0] module_1_io_addr; // @[memory.scala 156:26]
  wire [31:0] module_1_io_data; // @[memory.scala 156:26]
  wire [1:0] module_1_io_size; // @[memory.scala 156:26]
  wire  module_1_io_en; // @[memory.scala 156:26]
  wire [9:0] module_1_io_mem_addr; // @[memory.scala 156:26]
  wire [7:0] module_1_io_mem_data_0; // @[memory.scala 156:26]
  wire [7:0] module_1_io_mem_data_1; // @[memory.scala 156:26]
  wire [7:0] module_1_io_mem_data_2; // @[memory.scala 156:26]
  wire [7:0] module_1_io_mem_data_3; // @[memory.scala 156:26]
  wire  module_1_io_mem_masks_0; // @[memory.scala 156:26]
  wire  module_1_io_mem_masks_1; // @[memory.scala 156:26]
  wire  module_1_io_mem_masks_2; // @[memory.scala 156:26]
  wire  module_1_io_mem_masks_3; // @[memory.scala 156:26]
  wire [2:0] _io_core_ports_0_resp_bits_data_T_1 = io_core_ports_0_req_bits_typ - 3'h1; // @[memory.scala 60:24]
  wire [2:0] _io_core_ports_1_resp_bits_data_T_1 = io_core_ports_1_req_bits_typ - 3'h1; // @[memory.scala 60:24]
  wire [2:0] _io_debug_port_resp_bits_data_T_1 = io_debug_port_req_bits_typ - 3'h1; // @[memory.scala 60:24]
  MemReader_1stage MemReader_1stage_0 ( // @[memory.scala 120:26]
    .io_addr(io_core_ports_0_resp_bits_data_module_io_addr),
    .io_size(io_core_ports_0_resp_bits_data_module_io_size),
    .io_signed(io_core_ports_0_resp_bits_data_module_io_signed),
    .io_data(io_core_ports_0_resp_bits_data_module_io_data),
    .io_mem_addr(io_core_ports_0_resp_bits_data_module_io_mem_addr),
    .io_mem_data_0(io_core_ports_0_resp_bits_data_module_io_mem_data_0),
    .io_mem_data_1(io_core_ports_0_resp_bits_data_module_io_mem_data_1),
    .io_mem_data_2(io_core_ports_0_resp_bits_data_module_io_mem_data_2),
    .io_mem_data_3(io_core_ports_0_resp_bits_data_module_io_mem_data_3)
  );
  MemWriter_1stage MemWriter_1stage_0 ( // @[memory.scala 156:26]
    .io_addr(module__io_addr),
    .io_data(module__io_data),
    .io_size(module__io_size),
    .io_en(module__io_en),
    .io_mem_addr(module__io_mem_addr),
    .io_mem_data_0(module__io_mem_data_0),
    .io_mem_data_1(module__io_mem_data_1),
    .io_mem_data_2(module__io_mem_data_2),
    .io_mem_data_3(module__io_mem_data_3),
    .io_mem_masks_0(module__io_mem_masks_0),
    .io_mem_masks_1(module__io_mem_masks_1),
    .io_mem_masks_2(module__io_mem_masks_2),
    .io_mem_masks_3(module__io_mem_masks_3)
  );
  MemReader_1stage MemReader_1stage_1 ( // @[memory.scala 120:26]
    .io_addr(io_core_ports_1_resp_bits_data_module_io_addr),
    .io_size(io_core_ports_1_resp_bits_data_module_io_size),
    .io_signed(io_core_ports_1_resp_bits_data_module_io_signed),
    .io_data(io_core_ports_1_resp_bits_data_module_io_data),
    .io_mem_addr(io_core_ports_1_resp_bits_data_module_io_mem_addr),
    .io_mem_data_0(io_core_ports_1_resp_bits_data_module_io_mem_data_0),
    .io_mem_data_1(io_core_ports_1_resp_bits_data_module_io_mem_data_1),
    .io_mem_data_2(io_core_ports_1_resp_bits_data_module_io_mem_data_2),
    .io_mem_data_3(io_core_ports_1_resp_bits_data_module_io_mem_data_3)
  );
  MemReader_1stage MemReader_1stage_2 ( // @[memory.scala 120:26]
    .io_addr(io_debug_port_resp_bits_data_module_io_addr),
    .io_size(io_debug_port_resp_bits_data_module_io_size),
    .io_signed(io_debug_port_resp_bits_data_module_io_signed),
    .io_data(io_debug_port_resp_bits_data_module_io_data),
    .io_mem_addr(io_debug_port_resp_bits_data_module_io_mem_addr),
    .io_mem_data_0(io_debug_port_resp_bits_data_module_io_mem_data_0),
    .io_mem_data_1(io_debug_port_resp_bits_data_module_io_mem_data_1),
    .io_mem_data_2(io_debug_port_resp_bits_data_module_io_mem_data_2),
    .io_mem_data_3(io_debug_port_resp_bits_data_module_io_mem_data_3)
  );
  MemWriter_1stage MemWriter_1stage_1 ( // @[memory.scala 156:26]
    .io_addr(module_1_io_addr),
    .io_data(module_1_io_data),
    .io_size(module_1_io_size),
    .io_en(module_1_io_en),
    .io_mem_addr(module_1_io_mem_addr),
    .io_mem_data_0(module_1_io_mem_data_0),
    .io_mem_data_1(module_1_io_mem_data_1),
    .io_mem_data_2(module_1_io_mem_data_2),
    .io_mem_data_3(module_1_io_mem_data_3),
    .io_mem_masks_0(module_1_io_mem_masks_0),
    .io_mem_masks_1(module_1_io_mem_masks_1),
    .io_mem_masks_2(module_1_io_mem_masks_2),
    .io_mem_masks_3(module_1_io_mem_masks_3)
  );
  assign mem_0_io_core_ports_0_resp_bits_data_MPORT_en = 1'h1;
  assign mem_0_io_core_ports_0_resp_bits_data_MPORT_addr = io_core_ports_0_resp_bits_data_module_io_mem_addr;
  assign mem_0_io_core_ports_0_resp_bits_data_MPORT_data = mem_0_0[mem_0_io_core_ports_0_resp_bits_data_MPORT_addr]; // @[memory.scala 73:31]
  assign mem_0_io_core_ports_1_resp_bits_data_MPORT_en = 1'h1;
  assign mem_0_io_core_ports_1_resp_bits_data_MPORT_addr = io_core_ports_1_resp_bits_data_module_io_mem_addr;
  assign mem_0_io_core_ports_1_resp_bits_data_MPORT_data = mem_0_1[mem_0_io_core_ports_1_resp_bits_data_MPORT_addr]; // @[memory.scala 73:31]
  assign mem_0_io_debug_port_resp_bits_data_MPORT_en = 1'h1;
  assign mem_0_io_debug_port_resp_bits_data_MPORT_addr = io_debug_port_resp_bits_data_module_io_mem_addr;
  assign mem_0_io_debug_port_resp_bits_data_MPORT_data = mem_0_0[mem_0_io_debug_port_resp_bits_data_MPORT_addr]; // @[memory.scala 73:31]
  assign mem_0_MPORT_data = module__io_mem_data_0;
  assign mem_0_MPORT_addr = module__io_mem_addr;
  assign mem_0_MPORT_mask = module__io_mem_masks_0;
  assign mem_0_MPORT_en = io_core_ports_0_req_valid & io_core_ports_0_req_bits_fcn;
  assign mem_0_MPORT_1_data = module_1_io_mem_data_0;
  assign mem_0_MPORT_1_addr = module_1_io_mem_addr;
  assign mem_0_MPORT_1_mask = module_1_io_mem_masks_0;
  assign mem_0_MPORT_1_en = io_debug_port_req_valid & io_debug_port_req_bits_fcn;
  assign mem_1_io_core_ports_0_resp_bits_data_MPORT_en = 1'h1;
  assign mem_1_io_core_ports_0_resp_bits_data_MPORT_addr = io_core_ports_0_resp_bits_data_module_io_mem_addr;
  assign mem_1_io_core_ports_0_resp_bits_data_MPORT_data = mem_1_0[mem_1_io_core_ports_0_resp_bits_data_MPORT_addr]; // @[memory.scala 73:31]
  assign mem_1_io_core_ports_1_resp_bits_data_MPORT_en = 1'h1;
  assign mem_1_io_core_ports_1_resp_bits_data_MPORT_addr = io_core_ports_1_resp_bits_data_module_io_mem_addr;
  assign mem_1_io_core_ports_1_resp_bits_data_MPORT_data = mem_1_1[mem_1_io_core_ports_1_resp_bits_data_MPORT_addr]; // @[memory.scala 73:31]
  assign mem_1_io_debug_port_resp_bits_data_MPORT_en = 1'h1;
  assign mem_1_io_debug_port_resp_bits_data_MPORT_addr = io_debug_port_resp_bits_data_module_io_mem_addr;
  assign mem_1_io_debug_port_resp_bits_data_MPORT_data = mem_1_0[mem_1_io_debug_port_resp_bits_data_MPORT_addr]; // @[memory.scala 73:31]
  assign mem_1_MPORT_data = module__io_mem_data_1;
  assign mem_1_MPORT_addr = module__io_mem_addr;
  assign mem_1_MPORT_mask = module__io_mem_masks_1;
  assign mem_1_MPORT_en = io_core_ports_0_req_valid & io_core_ports_0_req_bits_fcn;
  assign mem_1_MPORT_1_data = module_1_io_mem_data_1;
  assign mem_1_MPORT_1_addr = module_1_io_mem_addr;
  assign mem_1_MPORT_1_mask = module_1_io_mem_masks_1;
  assign mem_1_MPORT_1_en = io_debug_port_req_valid & io_debug_port_req_bits_fcn;
  assign mem_2_io_core_ports_0_resp_bits_data_MPORT_en = 1'h1;
  assign mem_2_io_core_ports_0_resp_bits_data_MPORT_addr = io_core_ports_0_resp_bits_data_module_io_mem_addr;
  assign mem_2_io_core_ports_0_resp_bits_data_MPORT_data = mem_2_0[mem_2_io_core_ports_0_resp_bits_data_MPORT_addr]; // @[memory.scala 73:31]
  assign mem_2_io_core_ports_1_resp_bits_data_MPORT_en = 1'h1;
  assign mem_2_io_core_ports_1_resp_bits_data_MPORT_addr = io_core_ports_1_resp_bits_data_module_io_mem_addr;
  assign mem_2_io_core_ports_1_resp_bits_data_MPORT_data = mem_2_1[mem_2_io_core_ports_1_resp_bits_data_MPORT_addr]; // @[memory.scala 73:31]
  assign mem_2_io_debug_port_resp_bits_data_MPORT_en = 1'h1;
  assign mem_2_io_debug_port_resp_bits_data_MPORT_addr = io_debug_port_resp_bits_data_module_io_mem_addr;
  assign mem_2_io_debug_port_resp_bits_data_MPORT_data = mem_2_0[mem_2_io_debug_port_resp_bits_data_MPORT_addr]; // @[memory.scala 73:31]
  assign mem_2_MPORT_data = module__io_mem_data_2;
  assign mem_2_MPORT_addr = module__io_mem_addr;
  assign mem_2_MPORT_mask = module__io_mem_masks_2;
  assign mem_2_MPORT_en = io_core_ports_0_req_valid & io_core_ports_0_req_bits_fcn;
  assign mem_2_MPORT_1_data = module_1_io_mem_data_2;
  assign mem_2_MPORT_1_addr = module_1_io_mem_addr;
  assign mem_2_MPORT_1_mask = module_1_io_mem_masks_2;
  assign mem_2_MPORT_1_en = io_debug_port_req_valid & io_debug_port_req_bits_fcn;
  assign mem_3_io_core_ports_0_resp_bits_data_MPORT_en = 1'h1;
  assign mem_3_io_core_ports_0_resp_bits_data_MPORT_addr = io_core_ports_0_resp_bits_data_module_io_mem_addr;
  assign mem_3_io_core_ports_0_resp_bits_data_MPORT_data = mem_3_0[mem_3_io_core_ports_0_resp_bits_data_MPORT_addr]; // @[memory.scala 73:31]
  assign mem_3_io_core_ports_1_resp_bits_data_MPORT_en = 1'h1;
  assign mem_3_io_core_ports_1_resp_bits_data_MPORT_addr = io_core_ports_1_resp_bits_data_module_io_mem_addr;
  assign mem_3_io_core_ports_1_resp_bits_data_MPORT_data = mem_3_1[mem_3_io_core_ports_1_resp_bits_data_MPORT_addr]; // @[memory.scala 73:31]
  assign mem_3_io_debug_port_resp_bits_data_MPORT_en = 1'h1;
  assign mem_3_io_debug_port_resp_bits_data_MPORT_addr = io_debug_port_resp_bits_data_module_io_mem_addr;
  assign mem_3_io_debug_port_resp_bits_data_MPORT_data = mem_3_0[mem_3_io_debug_port_resp_bits_data_MPORT_addr]; // @[memory.scala 73:31]
  assign mem_3_MPORT_data = module__io_mem_data_3;
  assign mem_3_MPORT_addr = module__io_mem_addr;
  assign mem_3_MPORT_mask = module__io_mem_masks_3;
  assign mem_3_MPORT_en = io_core_ports_0_req_valid & io_core_ports_0_req_bits_fcn;
  assign mem_3_MPORT_1_data = module_1_io_mem_data_3;
  assign mem_3_MPORT_1_addr = module_1_io_mem_addr;
  assign mem_3_MPORT_1_mask = module_1_io_mem_masks_3;
  assign mem_3_MPORT_1_en = io_debug_port_req_valid & io_debug_port_req_bits_fcn;
  assign io_core_ports_0_resp_valid = io_core_ports_0_req_valid; // @[memory.scala 185:35]
  assign io_core_ports_0_resp_bits_data = io_core_ports_0_resp_bits_data_module_io_data; // @[memory.scala 194:40]
  assign io_core_ports_1_resp_valid = io_core_ports_1_req_valid; // @[memory.scala 185:35]
  assign io_core_ports_1_resp_bits_data = io_core_ports_1_resp_bits_data_module_io_data; // @[memory.scala 201:43]
  assign io_debug_port_resp_valid = io_debug_port_req_valid; // @[memory.scala 207:29]
  assign io_debug_port_resp_bits_data = io_debug_port_resp_bits_data_module_io_data; // @[memory.scala 211:33]
  assign io_core_ports_0_resp_bits_data_module_io_addr = io_core_ports_0_req_bits_addr[20:0]; // @[memory.scala 121:22]
  assign io_core_ports_0_resp_bits_data_module_io_size = _io_core_ports_0_resp_bits_data_T_1[1:0]; // @[memory.scala 60:30]
  assign io_core_ports_0_resp_bits_data_module_io_signed = ~_io_core_ports_0_resp_bits_data_T_1[2]; // @[memory.scala 61:21]
  assign io_core_ports_0_resp_bits_data_module_io_mem_data_0 = mem_0_io_core_ports_0_resp_bits_data_MPORT_data; // @[memory.scala 124:26]
  assign io_core_ports_0_resp_bits_data_module_io_mem_data_1 = mem_1_io_core_ports_0_resp_bits_data_MPORT_data; // @[memory.scala 124:26]
  assign io_core_ports_0_resp_bits_data_module_io_mem_data_2 = mem_2_io_core_ports_0_resp_bits_data_MPORT_data; // @[memory.scala 124:26]
  assign io_core_ports_0_resp_bits_data_module_io_mem_data_3 = mem_3_io_core_ports_0_resp_bits_data_MPORT_data; // @[memory.scala 124:26]
  assign module__io_addr = io_core_ports_0_req_bits_addr[20:0]; // @[memory.scala 157:22]
  assign module__io_data = io_core_ports_0_req_bits_data; // @[memory.scala 158:22]
  assign module__io_size = _io_core_ports_0_resp_bits_data_T_1[1:0]; // @[memory.scala 60:30]
  assign module__io_en = io_core_ports_0_req_valid & io_core_ports_0_req_bits_fcn; // @[memory.scala 193:51]
  assign io_core_ports_1_resp_bits_data_module_io_addr = io_core_ports_1_req_bits_addr[20:0]; // @[memory.scala 121:22]
  assign io_core_ports_1_resp_bits_data_module_io_size = _io_core_ports_1_resp_bits_data_T_1[1:0]; // @[memory.scala 60:30]
  assign io_core_ports_1_resp_bits_data_module_io_signed = ~_io_core_ports_1_resp_bits_data_T_1[2]; // @[memory.scala 61:21]
  assign io_core_ports_1_resp_bits_data_module_io_mem_data_0 = mem_0_io_core_ports_1_resp_bits_data_MPORT_data; // @[memory.scala 124:26]
  assign io_core_ports_1_resp_bits_data_module_io_mem_data_1 = mem_1_io_core_ports_1_resp_bits_data_MPORT_data; // @[memory.scala 124:26]
  assign io_core_ports_1_resp_bits_data_module_io_mem_data_2 = mem_2_io_core_ports_1_resp_bits_data_MPORT_data; // @[memory.scala 124:26]
  assign io_core_ports_1_resp_bits_data_module_io_mem_data_3 = mem_3_io_core_ports_1_resp_bits_data_MPORT_data; // @[memory.scala 124:26]
  assign io_debug_port_resp_bits_data_module_io_addr = io_debug_port_req_bits_addr[20:0]; // @[memory.scala 121:22]
  assign io_debug_port_resp_bits_data_module_io_size = _io_debug_port_resp_bits_data_T_1[1:0]; // @[memory.scala 60:30]
  assign io_debug_port_resp_bits_data_module_io_signed = ~_io_debug_port_resp_bits_data_T_1[2]; // @[memory.scala 61:21]
  assign io_debug_port_resp_bits_data_module_io_mem_data_0 = mem_0_io_debug_port_resp_bits_data_MPORT_data; // @[memory.scala 124:26]
  assign io_debug_port_resp_bits_data_module_io_mem_data_1 = mem_1_io_debug_port_resp_bits_data_MPORT_data; // @[memory.scala 124:26]
  assign io_debug_port_resp_bits_data_module_io_mem_data_2 = mem_2_io_debug_port_resp_bits_data_MPORT_data; // @[memory.scala 124:26]
  assign io_debug_port_resp_bits_data_module_io_mem_data_3 = mem_3_io_debug_port_resp_bits_data_MPORT_data; // @[memory.scala 124:26]
  assign module_1_io_addr = io_debug_port_req_bits_addr[20:0]; // @[memory.scala 157:22]
  assign module_1_io_data = io_debug_port_req_bits_data; // @[memory.scala 158:22]
  assign module_1_io_size = _io_debug_port_resp_bits_data_T_1[1:0]; // @[memory.scala 60:30]
  assign module_1_io_en = io_debug_port_req_valid & io_debug_port_req_bits_fcn; // @[memory.scala 210:49]
  always @(posedge clock) begin
    if (mem_0_MPORT_en & mem_0_MPORT_mask) begin
      mem_0_0[mem_0_MPORT_addr] <= mem_0_MPORT_data; // @[memory.scala 73:31]
    end
    if (mem_0_MPORT_1_en & mem_0_MPORT_1_mask) begin
      mem_0_0[mem_0_MPORT_1_addr] <= mem_0_MPORT_1_data; // @[memory.scala 73:31]
    end
    if (mem_1_MPORT_en & mem_1_MPORT_mask) begin
      mem_1_0[mem_1_MPORT_addr] <= mem_1_MPORT_data; // @[memory.scala 73:31]
    end
    if (mem_1_MPORT_1_en & mem_1_MPORT_1_mask) begin
      mem_1_0[mem_1_MPORT_1_addr] <= mem_1_MPORT_1_data; // @[memory.scala 73:31]
    end
    if (mem_2_MPORT_en & mem_2_MPORT_mask) begin
      mem_2_0[mem_2_MPORT_addr] <= mem_2_MPORT_data; // @[memory.scala 73:31]
    end
    if (mem_2_MPORT_1_en & mem_2_MPORT_1_mask) begin
      mem_2_0[mem_2_MPORT_1_addr] <= mem_2_MPORT_1_data; // @[memory.scala 73:31]
    end
    if (mem_3_MPORT_en & mem_3_MPORT_mask) begin
      mem_3_0[mem_3_MPORT_addr] <= mem_3_MPORT_data; // @[memory.scala 73:31]
    end
    if (mem_3_MPORT_1_en & mem_3_MPORT_1_mask) begin
      mem_3_0[mem_3_MPORT_1_addr] <= mem_3_MPORT_1_data; // @[memory.scala 73:31]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 524288; initvar = initvar+1)
    mem_0[initvar] = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 524288; initvar = initvar+1)
    mem_1[initvar] = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 524288; initvar = initvar+1)
    mem_2[initvar] = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 524288; initvar = initvar+1)
    mem_3[initvar] = _RAND_3[7:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
wire [8*(1024)-1:0] mem_0_1_flat_src;
assign mem_0_1_flat_src = {mem_0_1[0 + 0],mem_0_1[0 + 1],mem_0_1[0 + 2],mem_0_1[0 + 3],mem_0_1[0 + 4],mem_0_1[0 + 5],mem_0_1[0 + 6],mem_0_1[0 + 7],mem_0_1[0 + 8],mem_0_1[0 + 9],mem_0_1[0 + 10],mem_0_1[0 + 11],mem_0_1[0 + 12],mem_0_1[0 + 13],mem_0_1[0 + 14],mem_0_1[0 + 15],mem_0_1[0 + 16],mem_0_1[0 + 17],mem_0_1[0 + 18],mem_0_1[0 + 19],mem_0_1[0 + 20],mem_0_1[0 + 21],mem_0_1[0 + 22],mem_0_1[0 + 23],mem_0_1[0 + 24],mem_0_1[0 + 25],mem_0_1[0 + 26],mem_0_1[0 + 27],mem_0_1[0 + 28],mem_0_1[0 + 29],mem_0_1[0 + 30],mem_0_1[0 + 31],mem_0_1[0 + 32],mem_0_1[0 + 33],mem_0_1[0 + 34],mem_0_1[0 + 35],mem_0_1[0 + 36],mem_0_1[0 + 37],mem_0_1[0 + 38],mem_0_1[0 + 39],mem_0_1[0 + 40],mem_0_1[0 + 41],mem_0_1[0 + 42],mem_0_1[0 + 43],mem_0_1[0 + 44],mem_0_1[0 + 45],mem_0_1[0 + 46],mem_0_1[0 + 47],mem_0_1[0 + 48],mem_0_1[0 + 49],mem_0_1[0 + 50],mem_0_1[0 + 51],mem_0_1[0 + 52],mem_0_1[0 + 53],mem_0_1[0 + 54],mem_0_1[0 + 55],mem_0_1[0 + 56],mem_0_1[0 + 57],mem_0_1[0 + 58],mem_0_1[0 + 59],mem_0_1[0 + 60],mem_0_1[0 + 61],mem_0_1[0 + 62],mem_0_1[0 + 63],mem_0_1[0 + 64],mem_0_1[0 + 65],mem_0_1[0 + 66],mem_0_1[0 + 67],mem_0_1[0 + 68],mem_0_1[0 + 69],mem_0_1[0 + 70],mem_0_1[0 + 71],mem_0_1[0 + 72],mem_0_1[0 + 73],mem_0_1[0 + 74],mem_0_1[0 + 75],mem_0_1[0 + 76],mem_0_1[0 + 77],mem_0_1[0 + 78],mem_0_1[0 + 79],mem_0_1[0 + 80],mem_0_1[0 + 81],mem_0_1[0 + 82],mem_0_1[0 + 83],mem_0_1[0 + 84],mem_0_1[0 + 85],mem_0_1[0 + 86],mem_0_1[0 + 87],mem_0_1[0 + 88],mem_0_1[0 + 89],mem_0_1[0 + 90],mem_0_1[0 + 91],mem_0_1[0 + 92],mem_0_1[0 + 93],mem_0_1[0 + 94],mem_0_1[0 + 95],mem_0_1[0 + 96],mem_0_1[0 + 97],mem_0_1[0 + 98],mem_0_1[0 + 99],mem_0_1[0 + 100],mem_0_1[0 + 101],mem_0_1[0 + 102],mem_0_1[0 + 103],mem_0_1[0 + 104],mem_0_1[0 + 105],mem_0_1[0 + 106],mem_0_1[0 + 107],mem_0_1[0 + 108],mem_0_1[0 + 109],mem_0_1[0 + 110],mem_0_1[0 + 111],mem_0_1[0 + 112],mem_0_1[0 + 113],mem_0_1[0 + 114],mem_0_1[0 + 115],mem_0_1[0 + 116],mem_0_1[0 + 117],mem_0_1[0 + 118],mem_0_1[0 + 119],mem_0_1[0 + 120],mem_0_1[0 + 121],mem_0_1[0 + 122],mem_0_1[0 + 123],mem_0_1[0 + 124],mem_0_1[0 + 125],mem_0_1[0 + 126],mem_0_1[0 + 127],mem_0_1[0 + 128],mem_0_1[0 + 129],mem_0_1[0 + 130],mem_0_1[0 + 131],mem_0_1[0 + 132],mem_0_1[0 + 133],mem_0_1[0 + 134],mem_0_1[0 + 135],mem_0_1[0 + 136],mem_0_1[0 + 137],mem_0_1[0 + 138],mem_0_1[0 + 139],mem_0_1[0 + 140],mem_0_1[0 + 141],mem_0_1[0 + 142],mem_0_1[0 + 143],mem_0_1[0 + 144],mem_0_1[0 + 145],mem_0_1[0 + 146],mem_0_1[0 + 147],mem_0_1[0 + 148],mem_0_1[0 + 149],mem_0_1[0 + 150],mem_0_1[0 + 151],mem_0_1[0 + 152],mem_0_1[0 + 153],mem_0_1[0 + 154],mem_0_1[0 + 155],mem_0_1[0 + 156],mem_0_1[0 + 157],mem_0_1[0 + 158],mem_0_1[0 + 159],mem_0_1[0 + 160],mem_0_1[0 + 161],mem_0_1[0 + 162],mem_0_1[0 + 163],mem_0_1[0 + 164],mem_0_1[0 + 165],mem_0_1[0 + 166],mem_0_1[0 + 167],mem_0_1[0 + 168],mem_0_1[0 + 169],mem_0_1[0 + 170],mem_0_1[0 + 171],mem_0_1[0 + 172],mem_0_1[0 + 173],mem_0_1[0 + 174],mem_0_1[0 + 175],mem_0_1[0 + 176],mem_0_1[0 + 177],mem_0_1[0 + 178],mem_0_1[0 + 179],mem_0_1[0 + 180],mem_0_1[0 + 181],mem_0_1[0 + 182],mem_0_1[0 + 183],mem_0_1[0 + 184],mem_0_1[0 + 185],mem_0_1[0 + 186],mem_0_1[0 + 187],mem_0_1[0 + 188],mem_0_1[0 + 189],mem_0_1[0 + 190],mem_0_1[0 + 191],mem_0_1[0 + 192],mem_0_1[0 + 193],mem_0_1[0 + 194],mem_0_1[0 + 195],mem_0_1[0 + 196],mem_0_1[0 + 197],mem_0_1[0 + 198],mem_0_1[0 + 199],mem_0_1[0 + 200],mem_0_1[0 + 201],mem_0_1[0 + 202],mem_0_1[0 + 203],mem_0_1[0 + 204],mem_0_1[0 + 205],mem_0_1[0 + 206],mem_0_1[0 + 207],mem_0_1[0 + 208],mem_0_1[0 + 209],mem_0_1[0 + 210],mem_0_1[0 + 211],mem_0_1[0 + 212],mem_0_1[0 + 213],mem_0_1[0 + 214],mem_0_1[0 + 215],mem_0_1[0 + 216],mem_0_1[0 + 217],mem_0_1[0 + 218],mem_0_1[0 + 219],mem_0_1[0 + 220],mem_0_1[0 + 221],mem_0_1[0 + 222],mem_0_1[0 + 223],mem_0_1[0 + 224],mem_0_1[0 + 225],mem_0_1[0 + 226],mem_0_1[0 + 227],mem_0_1[0 + 228],mem_0_1[0 + 229],mem_0_1[0 + 230],mem_0_1[0 + 231],mem_0_1[0 + 232],mem_0_1[0 + 233],mem_0_1[0 + 234],mem_0_1[0 + 235],mem_0_1[0 + 236],mem_0_1[0 + 237],mem_0_1[0 + 238],mem_0_1[0 + 239],mem_0_1[0 + 240],mem_0_1[0 + 241],mem_0_1[0 + 242],mem_0_1[0 + 243],mem_0_1[0 + 244],mem_0_1[0 + 245],mem_0_1[0 + 246],mem_0_1[0 + 247],mem_0_1[0 + 248],mem_0_1[0 + 249],mem_0_1[0 + 250],mem_0_1[0 + 251],mem_0_1[0 + 252],mem_0_1[0 + 253],mem_0_1[0 + 254],mem_0_1[0 + 255],mem_0_1[0 + 256],mem_0_1[0 + 257],mem_0_1[0 + 258],mem_0_1[0 + 259],mem_0_1[0 + 260],mem_0_1[0 + 261],mem_0_1[0 + 262],mem_0_1[0 + 263],mem_0_1[0 + 264],mem_0_1[0 + 265],mem_0_1[0 + 266],mem_0_1[0 + 267],mem_0_1[0 + 268],mem_0_1[0 + 269],mem_0_1[0 + 270],mem_0_1[0 + 271],mem_0_1[0 + 272],mem_0_1[0 + 273],mem_0_1[0 + 274],mem_0_1[0 + 275],mem_0_1[0 + 276],mem_0_1[0 + 277],mem_0_1[0 + 278],mem_0_1[0 + 279],mem_0_1[0 + 280],mem_0_1[0 + 281],mem_0_1[0 + 282],mem_0_1[0 + 283],mem_0_1[0 + 284],mem_0_1[0 + 285],mem_0_1[0 + 286],mem_0_1[0 + 287],mem_0_1[0 + 288],mem_0_1[0 + 289],mem_0_1[0 + 290],mem_0_1[0 + 291],mem_0_1[0 + 292],mem_0_1[0 + 293],mem_0_1[0 + 294],mem_0_1[0 + 295],mem_0_1[0 + 296],mem_0_1[0 + 297],mem_0_1[0 + 298],mem_0_1[0 + 299],mem_0_1[0 + 300],mem_0_1[0 + 301],mem_0_1[0 + 302],mem_0_1[0 + 303],mem_0_1[0 + 304],mem_0_1[0 + 305],mem_0_1[0 + 306],mem_0_1[0 + 307],mem_0_1[0 + 308],mem_0_1[0 + 309],mem_0_1[0 + 310],mem_0_1[0 + 311],mem_0_1[0 + 312],mem_0_1[0 + 313],mem_0_1[0 + 314],mem_0_1[0 + 315],mem_0_1[0 + 316],mem_0_1[0 + 317],mem_0_1[0 + 318],mem_0_1[0 + 319],mem_0_1[0 + 320],mem_0_1[0 + 321],mem_0_1[0 + 322],mem_0_1[0 + 323],mem_0_1[0 + 324],mem_0_1[0 + 325],mem_0_1[0 + 326],mem_0_1[0 + 327],mem_0_1[0 + 328],mem_0_1[0 + 329],mem_0_1[0 + 330],mem_0_1[0 + 331],mem_0_1[0 + 332],mem_0_1[0 + 333],mem_0_1[0 + 334],mem_0_1[0 + 335],mem_0_1[0 + 336],mem_0_1[0 + 337],mem_0_1[0 + 338],mem_0_1[0 + 339],mem_0_1[0 + 340],mem_0_1[0 + 341],mem_0_1[0 + 342],mem_0_1[0 + 343],mem_0_1[0 + 344],mem_0_1[0 + 345],mem_0_1[0 + 346],mem_0_1[0 + 347],mem_0_1[0 + 348],mem_0_1[0 + 349],mem_0_1[0 + 350],mem_0_1[0 + 351],mem_0_1[0 + 352],mem_0_1[0 + 353],mem_0_1[0 + 354],mem_0_1[0 + 355],mem_0_1[0 + 356],mem_0_1[0 + 357],mem_0_1[0 + 358],mem_0_1[0 + 359],mem_0_1[0 + 360],mem_0_1[0 + 361],mem_0_1[0 + 362],mem_0_1[0 + 363],mem_0_1[0 + 364],mem_0_1[0 + 365],mem_0_1[0 + 366],mem_0_1[0 + 367],mem_0_1[0 + 368],mem_0_1[0 + 369],mem_0_1[0 + 370],mem_0_1[0 + 371],mem_0_1[0 + 372],mem_0_1[0 + 373],mem_0_1[0 + 374],mem_0_1[0 + 375],mem_0_1[0 + 376],mem_0_1[0 + 377],mem_0_1[0 + 378],mem_0_1[0 + 379],mem_0_1[0 + 380],mem_0_1[0 + 381],mem_0_1[0 + 382],mem_0_1[0 + 383],mem_0_1[0 + 384],mem_0_1[0 + 385],mem_0_1[0 + 386],mem_0_1[0 + 387],mem_0_1[0 + 388],mem_0_1[0 + 389],mem_0_1[0 + 390],mem_0_1[0 + 391],mem_0_1[0 + 392],mem_0_1[0 + 393],mem_0_1[0 + 394],mem_0_1[0 + 395],mem_0_1[0 + 396],mem_0_1[0 + 397],mem_0_1[0 + 398],mem_0_1[0 + 399],mem_0_1[0 + 400],mem_0_1[0 + 401],mem_0_1[0 + 402],mem_0_1[0 + 403],mem_0_1[0 + 404],mem_0_1[0 + 405],mem_0_1[0 + 406],mem_0_1[0 + 407],mem_0_1[0 + 408],mem_0_1[0 + 409],mem_0_1[0 + 410],mem_0_1[0 + 411],mem_0_1[0 + 412],mem_0_1[0 + 413],mem_0_1[0 + 414],mem_0_1[0 + 415],mem_0_1[0 + 416],mem_0_1[0 + 417],mem_0_1[0 + 418],mem_0_1[0 + 419],mem_0_1[0 + 420],mem_0_1[0 + 421],mem_0_1[0 + 422],mem_0_1[0 + 423],mem_0_1[0 + 424],mem_0_1[0 + 425],mem_0_1[0 + 426],mem_0_1[0 + 427],mem_0_1[0 + 428],mem_0_1[0 + 429],mem_0_1[0 + 430],mem_0_1[0 + 431],mem_0_1[0 + 432],mem_0_1[0 + 433],mem_0_1[0 + 434],mem_0_1[0 + 435],mem_0_1[0 + 436],mem_0_1[0 + 437],mem_0_1[0 + 438],mem_0_1[0 + 439],mem_0_1[0 + 440],mem_0_1[0 + 441],mem_0_1[0 + 442],mem_0_1[0 + 443],mem_0_1[0 + 444],mem_0_1[0 + 445],mem_0_1[0 + 446],mem_0_1[0 + 447],mem_0_1[0 + 448],mem_0_1[0 + 449],mem_0_1[0 + 450],mem_0_1[0 + 451],mem_0_1[0 + 452],mem_0_1[0 + 453],mem_0_1[0 + 454],mem_0_1[0 + 455],mem_0_1[0 + 456],mem_0_1[0 + 457],mem_0_1[0 + 458],mem_0_1[0 + 459],mem_0_1[0 + 460],mem_0_1[0 + 461],mem_0_1[0 + 462],mem_0_1[0 + 463],mem_0_1[0 + 464],mem_0_1[0 + 465],mem_0_1[0 + 466],mem_0_1[0 + 467],mem_0_1[0 + 468],mem_0_1[0 + 469],mem_0_1[0 + 470],mem_0_1[0 + 471],mem_0_1[0 + 472],mem_0_1[0 + 473],mem_0_1[0 + 474],mem_0_1[0 + 475],mem_0_1[0 + 476],mem_0_1[0 + 477],mem_0_1[0 + 478],mem_0_1[0 + 479],mem_0_1[0 + 480],mem_0_1[0 + 481],mem_0_1[0 + 482],mem_0_1[0 + 483],mem_0_1[0 + 484],mem_0_1[0 + 485],mem_0_1[0 + 486],mem_0_1[0 + 487],mem_0_1[0 + 488],mem_0_1[0 + 489],mem_0_1[0 + 490],mem_0_1[0 + 491],mem_0_1[0 + 492],mem_0_1[0 + 493],mem_0_1[0 + 494],mem_0_1[0 + 495],mem_0_1[0 + 496],mem_0_1[0 + 497],mem_0_1[0 + 498],mem_0_1[0 + 499],mem_0_1[0 + 500],mem_0_1[0 + 501],mem_0_1[0 + 502],mem_0_1[0 + 503],mem_0_1[0 + 504],mem_0_1[0 + 505],mem_0_1[0 + 506],mem_0_1[0 + 507],mem_0_1[0 + 508],mem_0_1[0 + 509],mem_0_1[0 + 510],mem_0_1[0 + 511],mem_0_1[0 + 512],mem_0_1[0 + 513],mem_0_1[0 + 514],mem_0_1[0 + 515],mem_0_1[0 + 516],mem_0_1[0 + 517],mem_0_1[0 + 518],mem_0_1[0 + 519],mem_0_1[0 + 520],mem_0_1[0 + 521],mem_0_1[0 + 522],mem_0_1[0 + 523],mem_0_1[0 + 524],mem_0_1[0 + 525],mem_0_1[0 + 526],mem_0_1[0 + 527],mem_0_1[0 + 528],mem_0_1[0 + 529],mem_0_1[0 + 530],mem_0_1[0 + 531],mem_0_1[0 + 532],mem_0_1[0 + 533],mem_0_1[0 + 534],mem_0_1[0 + 535],mem_0_1[0 + 536],mem_0_1[0 + 537],mem_0_1[0 + 538],mem_0_1[0 + 539],mem_0_1[0 + 540],mem_0_1[0 + 541],mem_0_1[0 + 542],mem_0_1[0 + 543],mem_0_1[0 + 544],mem_0_1[0 + 545],mem_0_1[0 + 546],mem_0_1[0 + 547],mem_0_1[0 + 548],mem_0_1[0 + 549],mem_0_1[0 + 550],mem_0_1[0 + 551],mem_0_1[0 + 552],mem_0_1[0 + 553],mem_0_1[0 + 554],mem_0_1[0 + 555],mem_0_1[0 + 556],mem_0_1[0 + 557],mem_0_1[0 + 558],mem_0_1[0 + 559],mem_0_1[0 + 560],mem_0_1[0 + 561],mem_0_1[0 + 562],mem_0_1[0 + 563],mem_0_1[0 + 564],mem_0_1[0 + 565],mem_0_1[0 + 566],mem_0_1[0 + 567],mem_0_1[0 + 568],mem_0_1[0 + 569],mem_0_1[0 + 570],mem_0_1[0 + 571],mem_0_1[0 + 572],mem_0_1[0 + 573],mem_0_1[0 + 574],mem_0_1[0 + 575],mem_0_1[0 + 576],mem_0_1[0 + 577],mem_0_1[0 + 578],mem_0_1[0 + 579],mem_0_1[0 + 580],mem_0_1[0 + 581],mem_0_1[0 + 582],mem_0_1[0 + 583],mem_0_1[0 + 584],mem_0_1[0 + 585],mem_0_1[0 + 586],mem_0_1[0 + 587],mem_0_1[0 + 588],mem_0_1[0 + 589],mem_0_1[0 + 590],mem_0_1[0 + 591],mem_0_1[0 + 592],mem_0_1[0 + 593],mem_0_1[0 + 594],mem_0_1[0 + 595],mem_0_1[0 + 596],mem_0_1[0 + 597],mem_0_1[0 + 598],mem_0_1[0 + 599],mem_0_1[0 + 600],mem_0_1[0 + 601],mem_0_1[0 + 602],mem_0_1[0 + 603],mem_0_1[0 + 604],mem_0_1[0 + 605],mem_0_1[0 + 606],mem_0_1[0 + 607],mem_0_1[0 + 608],mem_0_1[0 + 609],mem_0_1[0 + 610],mem_0_1[0 + 611],mem_0_1[0 + 612],mem_0_1[0 + 613],mem_0_1[0 + 614],mem_0_1[0 + 615],mem_0_1[0 + 616],mem_0_1[0 + 617],mem_0_1[0 + 618],mem_0_1[0 + 619],mem_0_1[0 + 620],mem_0_1[0 + 621],mem_0_1[0 + 622],mem_0_1[0 + 623],mem_0_1[0 + 624],mem_0_1[0 + 625],mem_0_1[0 + 626],mem_0_1[0 + 627],mem_0_1[0 + 628],mem_0_1[0 + 629],mem_0_1[0 + 630],mem_0_1[0 + 631],mem_0_1[0 + 632],mem_0_1[0 + 633],mem_0_1[0 + 634],mem_0_1[0 + 635],mem_0_1[0 + 636],mem_0_1[0 + 637],mem_0_1[0 + 638],mem_0_1[0 + 639],mem_0_1[0 + 640],mem_0_1[0 + 641],mem_0_1[0 + 642],mem_0_1[0 + 643],mem_0_1[0 + 644],mem_0_1[0 + 645],mem_0_1[0 + 646],mem_0_1[0 + 647],mem_0_1[0 + 648],mem_0_1[0 + 649],mem_0_1[0 + 650],mem_0_1[0 + 651],mem_0_1[0 + 652],mem_0_1[0 + 653],mem_0_1[0 + 654],mem_0_1[0 + 655],mem_0_1[0 + 656],mem_0_1[0 + 657],mem_0_1[0 + 658],mem_0_1[0 + 659],mem_0_1[0 + 660],mem_0_1[0 + 661],mem_0_1[0 + 662],mem_0_1[0 + 663],mem_0_1[0 + 664],mem_0_1[0 + 665],mem_0_1[0 + 666],mem_0_1[0 + 667],mem_0_1[0 + 668],mem_0_1[0 + 669],mem_0_1[0 + 670],mem_0_1[0 + 671],mem_0_1[0 + 672],mem_0_1[0 + 673],mem_0_1[0 + 674],mem_0_1[0 + 675],mem_0_1[0 + 676],mem_0_1[0 + 677],mem_0_1[0 + 678],mem_0_1[0 + 679],mem_0_1[0 + 680],mem_0_1[0 + 681],mem_0_1[0 + 682],mem_0_1[0 + 683],mem_0_1[0 + 684],mem_0_1[0 + 685],mem_0_1[0 + 686],mem_0_1[0 + 687],mem_0_1[0 + 688],mem_0_1[0 + 689],mem_0_1[0 + 690],mem_0_1[0 + 691],mem_0_1[0 + 692],mem_0_1[0 + 693],mem_0_1[0 + 694],mem_0_1[0 + 695],mem_0_1[0 + 696],mem_0_1[0 + 697],mem_0_1[0 + 698],mem_0_1[0 + 699],mem_0_1[0 + 700],mem_0_1[0 + 701],mem_0_1[0 + 702],mem_0_1[0 + 703],mem_0_1[0 + 704],mem_0_1[0 + 705],mem_0_1[0 + 706],mem_0_1[0 + 707],mem_0_1[0 + 708],mem_0_1[0 + 709],mem_0_1[0 + 710],mem_0_1[0 + 711],mem_0_1[0 + 712],mem_0_1[0 + 713],mem_0_1[0 + 714],mem_0_1[0 + 715],mem_0_1[0 + 716],mem_0_1[0 + 717],mem_0_1[0 + 718],mem_0_1[0 + 719],mem_0_1[0 + 720],mem_0_1[0 + 721],mem_0_1[0 + 722],mem_0_1[0 + 723],mem_0_1[0 + 724],mem_0_1[0 + 725],mem_0_1[0 + 726],mem_0_1[0 + 727],mem_0_1[0 + 728],mem_0_1[0 + 729],mem_0_1[0 + 730],mem_0_1[0 + 731],mem_0_1[0 + 732],mem_0_1[0 + 733],mem_0_1[0 + 734],mem_0_1[0 + 735],mem_0_1[0 + 736],mem_0_1[0 + 737],mem_0_1[0 + 738],mem_0_1[0 + 739],mem_0_1[0 + 740],mem_0_1[0 + 741],mem_0_1[0 + 742],mem_0_1[0 + 743],mem_0_1[0 + 744],mem_0_1[0 + 745],mem_0_1[0 + 746],mem_0_1[0 + 747],mem_0_1[0 + 748],mem_0_1[0 + 749],mem_0_1[0 + 750],mem_0_1[0 + 751],mem_0_1[0 + 752],mem_0_1[0 + 753],mem_0_1[0 + 754],mem_0_1[0 + 755],mem_0_1[0 + 756],mem_0_1[0 + 757],mem_0_1[0 + 758],mem_0_1[0 + 759],mem_0_1[0 + 760],mem_0_1[0 + 761],mem_0_1[0 + 762],mem_0_1[0 + 763],mem_0_1[0 + 764],mem_0_1[0 + 765],mem_0_1[0 + 766],mem_0_1[0 + 767],mem_0_1[0 + 768],mem_0_1[0 + 769],mem_0_1[0 + 770],mem_0_1[0 + 771],mem_0_1[0 + 772],mem_0_1[0 + 773],mem_0_1[0 + 774],mem_0_1[0 + 775],mem_0_1[0 + 776],mem_0_1[0 + 777],mem_0_1[0 + 778],mem_0_1[0 + 779],mem_0_1[0 + 780],mem_0_1[0 + 781],mem_0_1[0 + 782],mem_0_1[0 + 783],mem_0_1[0 + 784],mem_0_1[0 + 785],mem_0_1[0 + 786],mem_0_1[0 + 787],mem_0_1[0 + 788],mem_0_1[0 + 789],mem_0_1[0 + 790],mem_0_1[0 + 791],mem_0_1[0 + 792],mem_0_1[0 + 793],mem_0_1[0 + 794],mem_0_1[0 + 795],mem_0_1[0 + 796],mem_0_1[0 + 797],mem_0_1[0 + 798],mem_0_1[0 + 799],mem_0_1[0 + 800],mem_0_1[0 + 801],mem_0_1[0 + 802],mem_0_1[0 + 803],mem_0_1[0 + 804],mem_0_1[0 + 805],mem_0_1[0 + 806],mem_0_1[0 + 807],mem_0_1[0 + 808],mem_0_1[0 + 809],mem_0_1[0 + 810],mem_0_1[0 + 811],mem_0_1[0 + 812],mem_0_1[0 + 813],mem_0_1[0 + 814],mem_0_1[0 + 815],mem_0_1[0 + 816],mem_0_1[0 + 817],mem_0_1[0 + 818],mem_0_1[0 + 819],mem_0_1[0 + 820],mem_0_1[0 + 821],mem_0_1[0 + 822],mem_0_1[0 + 823],mem_0_1[0 + 824],mem_0_1[0 + 825],mem_0_1[0 + 826],mem_0_1[0 + 827],mem_0_1[0 + 828],mem_0_1[0 + 829],mem_0_1[0 + 830],mem_0_1[0 + 831],mem_0_1[0 + 832],mem_0_1[0 + 833],mem_0_1[0 + 834],mem_0_1[0 + 835],mem_0_1[0 + 836],mem_0_1[0 + 837],mem_0_1[0 + 838],mem_0_1[0 + 839],mem_0_1[0 + 840],mem_0_1[0 + 841],mem_0_1[0 + 842],mem_0_1[0 + 843],mem_0_1[0 + 844],mem_0_1[0 + 845],mem_0_1[0 + 846],mem_0_1[0 + 847],mem_0_1[0 + 848],mem_0_1[0 + 849],mem_0_1[0 + 850],mem_0_1[0 + 851],mem_0_1[0 + 852],mem_0_1[0 + 853],mem_0_1[0 + 854],mem_0_1[0 + 855],mem_0_1[0 + 856],mem_0_1[0 + 857],mem_0_1[0 + 858],mem_0_1[0 + 859],mem_0_1[0 + 860],mem_0_1[0 + 861],mem_0_1[0 + 862],mem_0_1[0 + 863],mem_0_1[0 + 864],mem_0_1[0 + 865],mem_0_1[0 + 866],mem_0_1[0 + 867],mem_0_1[0 + 868],mem_0_1[0 + 869],mem_0_1[0 + 870],mem_0_1[0 + 871],mem_0_1[0 + 872],mem_0_1[0 + 873],mem_0_1[0 + 874],mem_0_1[0 + 875],mem_0_1[0 + 876],mem_0_1[0 + 877],mem_0_1[0 + 878],mem_0_1[0 + 879],mem_0_1[0 + 880],mem_0_1[0 + 881],mem_0_1[0 + 882],mem_0_1[0 + 883],mem_0_1[0 + 884],mem_0_1[0 + 885],mem_0_1[0 + 886],mem_0_1[0 + 887],mem_0_1[0 + 888],mem_0_1[0 + 889],mem_0_1[0 + 890],mem_0_1[0 + 891],mem_0_1[0 + 892],mem_0_1[0 + 893],mem_0_1[0 + 894],mem_0_1[0 + 895],mem_0_1[0 + 896],mem_0_1[0 + 897],mem_0_1[0 + 898],mem_0_1[0 + 899],mem_0_1[0 + 900],mem_0_1[0 + 901],mem_0_1[0 + 902],mem_0_1[0 + 903],mem_0_1[0 + 904],mem_0_1[0 + 905],mem_0_1[0 + 906],mem_0_1[0 + 907],mem_0_1[0 + 908],mem_0_1[0 + 909],mem_0_1[0 + 910],mem_0_1[0 + 911],mem_0_1[0 + 912],mem_0_1[0 + 913],mem_0_1[0 + 914],mem_0_1[0 + 915],mem_0_1[0 + 916],mem_0_1[0 + 917],mem_0_1[0 + 918],mem_0_1[0 + 919],mem_0_1[0 + 920],mem_0_1[0 + 921],mem_0_1[0 + 922],mem_0_1[0 + 923],mem_0_1[0 + 924],mem_0_1[0 + 925],mem_0_1[0 + 926],mem_0_1[0 + 927],mem_0_1[0 + 928],mem_0_1[0 + 929],mem_0_1[0 + 930],mem_0_1[0 + 931],mem_0_1[0 + 932],mem_0_1[0 + 933],mem_0_1[0 + 934],mem_0_1[0 + 935],mem_0_1[0 + 936],mem_0_1[0 + 937],mem_0_1[0 + 938],mem_0_1[0 + 939],mem_0_1[0 + 940],mem_0_1[0 + 941],mem_0_1[0 + 942],mem_0_1[0 + 943],mem_0_1[0 + 944],mem_0_1[0 + 945],mem_0_1[0 + 946],mem_0_1[0 + 947],mem_0_1[0 + 948],mem_0_1[0 + 949],mem_0_1[0 + 950],mem_0_1[0 + 951],mem_0_1[0 + 952],mem_0_1[0 + 953],mem_0_1[0 + 954],mem_0_1[0 + 955],mem_0_1[0 + 956],mem_0_1[0 + 957],mem_0_1[0 + 958],mem_0_1[0 + 959],mem_0_1[0 + 960],mem_0_1[0 + 961],mem_0_1[0 + 962],mem_0_1[0 + 963],mem_0_1[0 + 964],mem_0_1[0 + 965],mem_0_1[0 + 966],mem_0_1[0 + 967],mem_0_1[0 + 968],mem_0_1[0 + 969],mem_0_1[0 + 970],mem_0_1[0 + 971],mem_0_1[0 + 972],mem_0_1[0 + 973],mem_0_1[0 + 974],mem_0_1[0 + 975],mem_0_1[0 + 976],mem_0_1[0 + 977],mem_0_1[0 + 978],mem_0_1[0 + 979],mem_0_1[0 + 980],mem_0_1[0 + 981],mem_0_1[0 + 982],mem_0_1[0 + 983],mem_0_1[0 + 984],mem_0_1[0 + 985],mem_0_1[0 + 986],mem_0_1[0 + 987],mem_0_1[0 + 988],mem_0_1[0 + 989],mem_0_1[0 + 990],mem_0_1[0 + 991],mem_0_1[0 + 992],mem_0_1[0 + 993],mem_0_1[0 + 994],mem_0_1[0 + 995],mem_0_1[0 + 996],mem_0_1[0 + 997],mem_0_1[0 + 998],mem_0_1[0 + 999],mem_0_1[0 + 1000],mem_0_1[0 + 1001],mem_0_1[0 + 1002],mem_0_1[0 + 1003],mem_0_1[0 + 1004],mem_0_1[0 + 1005],mem_0_1[0 + 1006],mem_0_1[0 + 1007],mem_0_1[0 + 1008],mem_0_1[0 + 1009],mem_0_1[0 + 1010],mem_0_1[0 + 1011],mem_0_1[0 + 1012],mem_0_1[0 + 1013],mem_0_1[0 + 1014],mem_0_1[0 + 1015],mem_0_1[0 + 1016],mem_0_1[0 + 1017],mem_0_1[0 + 1018],mem_0_1[0 + 1019],mem_0_1[0 + 1020],mem_0_1[0 + 1021],mem_0_1[0 + 1022],mem_0_1[0 + 1024 - 1] };
wire [8*(1024)-1:0] mem_1_1_flat_src;
assign mem_1_1_flat_src = {mem_1_1[0 + 0],mem_1_1[0 + 1],mem_1_1[0 + 2],mem_1_1[0 + 3],mem_1_1[0 + 4],mem_1_1[0 + 5],mem_1_1[0 + 6],mem_1_1[0 + 7],mem_1_1[0 + 8],mem_1_1[0 + 9],mem_1_1[0 + 10],mem_1_1[0 + 11],mem_1_1[0 + 12],mem_1_1[0 + 13],mem_1_1[0 + 14],mem_1_1[0 + 15],mem_1_1[0 + 16],mem_1_1[0 + 17],mem_1_1[0 + 18],mem_1_1[0 + 19],mem_1_1[0 + 20],mem_1_1[0 + 21],mem_1_1[0 + 22],mem_1_1[0 + 23],mem_1_1[0 + 24],mem_1_1[0 + 25],mem_1_1[0 + 26],mem_1_1[0 + 27],mem_1_1[0 + 28],mem_1_1[0 + 29],mem_1_1[0 + 30],mem_1_1[0 + 31],mem_1_1[0 + 32],mem_1_1[0 + 33],mem_1_1[0 + 34],mem_1_1[0 + 35],mem_1_1[0 + 36],mem_1_1[0 + 37],mem_1_1[0 + 38],mem_1_1[0 + 39],mem_1_1[0 + 40],mem_1_1[0 + 41],mem_1_1[0 + 42],mem_1_1[0 + 43],mem_1_1[0 + 44],mem_1_1[0 + 45],mem_1_1[0 + 46],mem_1_1[0 + 47],mem_1_1[0 + 48],mem_1_1[0 + 49],mem_1_1[0 + 50],mem_1_1[0 + 51],mem_1_1[0 + 52],mem_1_1[0 + 53],mem_1_1[0 + 54],mem_1_1[0 + 55],mem_1_1[0 + 56],mem_1_1[0 + 57],mem_1_1[0 + 58],mem_1_1[0 + 59],mem_1_1[0 + 60],mem_1_1[0 + 61],mem_1_1[0 + 62],mem_1_1[0 + 63],mem_1_1[0 + 64],mem_1_1[0 + 65],mem_1_1[0 + 66],mem_1_1[0 + 67],mem_1_1[0 + 68],mem_1_1[0 + 69],mem_1_1[0 + 70],mem_1_1[0 + 71],mem_1_1[0 + 72],mem_1_1[0 + 73],mem_1_1[0 + 74],mem_1_1[0 + 75],mem_1_1[0 + 76],mem_1_1[0 + 77],mem_1_1[0 + 78],mem_1_1[0 + 79],mem_1_1[0 + 80],mem_1_1[0 + 81],mem_1_1[0 + 82],mem_1_1[0 + 83],mem_1_1[0 + 84],mem_1_1[0 + 85],mem_1_1[0 + 86],mem_1_1[0 + 87],mem_1_1[0 + 88],mem_1_1[0 + 89],mem_1_1[0 + 90],mem_1_1[0 + 91],mem_1_1[0 + 92],mem_1_1[0 + 93],mem_1_1[0 + 94],mem_1_1[0 + 95],mem_1_1[0 + 96],mem_1_1[0 + 97],mem_1_1[0 + 98],mem_1_1[0 + 99],mem_1_1[0 + 100],mem_1_1[0 + 101],mem_1_1[0 + 102],mem_1_1[0 + 103],mem_1_1[0 + 104],mem_1_1[0 + 105],mem_1_1[0 + 106],mem_1_1[0 + 107],mem_1_1[0 + 108],mem_1_1[0 + 109],mem_1_1[0 + 110],mem_1_1[0 + 111],mem_1_1[0 + 112],mem_1_1[0 + 113],mem_1_1[0 + 114],mem_1_1[0 + 115],mem_1_1[0 + 116],mem_1_1[0 + 117],mem_1_1[0 + 118],mem_1_1[0 + 119],mem_1_1[0 + 120],mem_1_1[0 + 121],mem_1_1[0 + 122],mem_1_1[0 + 123],mem_1_1[0 + 124],mem_1_1[0 + 125],mem_1_1[0 + 126],mem_1_1[0 + 127],mem_1_1[0 + 128],mem_1_1[0 + 129],mem_1_1[0 + 130],mem_1_1[0 + 131],mem_1_1[0 + 132],mem_1_1[0 + 133],mem_1_1[0 + 134],mem_1_1[0 + 135],mem_1_1[0 + 136],mem_1_1[0 + 137],mem_1_1[0 + 138],mem_1_1[0 + 139],mem_1_1[0 + 140],mem_1_1[0 + 141],mem_1_1[0 + 142],mem_1_1[0 + 143],mem_1_1[0 + 144],mem_1_1[0 + 145],mem_1_1[0 + 146],mem_1_1[0 + 147],mem_1_1[0 + 148],mem_1_1[0 + 149],mem_1_1[0 + 150],mem_1_1[0 + 151],mem_1_1[0 + 152],mem_1_1[0 + 153],mem_1_1[0 + 154],mem_1_1[0 + 155],mem_1_1[0 + 156],mem_1_1[0 + 157],mem_1_1[0 + 158],mem_1_1[0 + 159],mem_1_1[0 + 160],mem_1_1[0 + 161],mem_1_1[0 + 162],mem_1_1[0 + 163],mem_1_1[0 + 164],mem_1_1[0 + 165],mem_1_1[0 + 166],mem_1_1[0 + 167],mem_1_1[0 + 168],mem_1_1[0 + 169],mem_1_1[0 + 170],mem_1_1[0 + 171],mem_1_1[0 + 172],mem_1_1[0 + 173],mem_1_1[0 + 174],mem_1_1[0 + 175],mem_1_1[0 + 176],mem_1_1[0 + 177],mem_1_1[0 + 178],mem_1_1[0 + 179],mem_1_1[0 + 180],mem_1_1[0 + 181],mem_1_1[0 + 182],mem_1_1[0 + 183],mem_1_1[0 + 184],mem_1_1[0 + 185],mem_1_1[0 + 186],mem_1_1[0 + 187],mem_1_1[0 + 188],mem_1_1[0 + 189],mem_1_1[0 + 190],mem_1_1[0 + 191],mem_1_1[0 + 192],mem_1_1[0 + 193],mem_1_1[0 + 194],mem_1_1[0 + 195],mem_1_1[0 + 196],mem_1_1[0 + 197],mem_1_1[0 + 198],mem_1_1[0 + 199],mem_1_1[0 + 200],mem_1_1[0 + 201],mem_1_1[0 + 202],mem_1_1[0 + 203],mem_1_1[0 + 204],mem_1_1[0 + 205],mem_1_1[0 + 206],mem_1_1[0 + 207],mem_1_1[0 + 208],mem_1_1[0 + 209],mem_1_1[0 + 210],mem_1_1[0 + 211],mem_1_1[0 + 212],mem_1_1[0 + 213],mem_1_1[0 + 214],mem_1_1[0 + 215],mem_1_1[0 + 216],mem_1_1[0 + 217],mem_1_1[0 + 218],mem_1_1[0 + 219],mem_1_1[0 + 220],mem_1_1[0 + 221],mem_1_1[0 + 222],mem_1_1[0 + 223],mem_1_1[0 + 224],mem_1_1[0 + 225],mem_1_1[0 + 226],mem_1_1[0 + 227],mem_1_1[0 + 228],mem_1_1[0 + 229],mem_1_1[0 + 230],mem_1_1[0 + 231],mem_1_1[0 + 232],mem_1_1[0 + 233],mem_1_1[0 + 234],mem_1_1[0 + 235],mem_1_1[0 + 236],mem_1_1[0 + 237],mem_1_1[0 + 238],mem_1_1[0 + 239],mem_1_1[0 + 240],mem_1_1[0 + 241],mem_1_1[0 + 242],mem_1_1[0 + 243],mem_1_1[0 + 244],mem_1_1[0 + 245],mem_1_1[0 + 246],mem_1_1[0 + 247],mem_1_1[0 + 248],mem_1_1[0 + 249],mem_1_1[0 + 250],mem_1_1[0 + 251],mem_1_1[0 + 252],mem_1_1[0 + 253],mem_1_1[0 + 254],mem_1_1[0 + 255],mem_1_1[0 + 256],mem_1_1[0 + 257],mem_1_1[0 + 258],mem_1_1[0 + 259],mem_1_1[0 + 260],mem_1_1[0 + 261],mem_1_1[0 + 262],mem_1_1[0 + 263],mem_1_1[0 + 264],mem_1_1[0 + 265],mem_1_1[0 + 266],mem_1_1[0 + 267],mem_1_1[0 + 268],mem_1_1[0 + 269],mem_1_1[0 + 270],mem_1_1[0 + 271],mem_1_1[0 + 272],mem_1_1[0 + 273],mem_1_1[0 + 274],mem_1_1[0 + 275],mem_1_1[0 + 276],mem_1_1[0 + 277],mem_1_1[0 + 278],mem_1_1[0 + 279],mem_1_1[0 + 280],mem_1_1[0 + 281],mem_1_1[0 + 282],mem_1_1[0 + 283],mem_1_1[0 + 284],mem_1_1[0 + 285],mem_1_1[0 + 286],mem_1_1[0 + 287],mem_1_1[0 + 288],mem_1_1[0 + 289],mem_1_1[0 + 290],mem_1_1[0 + 291],mem_1_1[0 + 292],mem_1_1[0 + 293],mem_1_1[0 + 294],mem_1_1[0 + 295],mem_1_1[0 + 296],mem_1_1[0 + 297],mem_1_1[0 + 298],mem_1_1[0 + 299],mem_1_1[0 + 300],mem_1_1[0 + 301],mem_1_1[0 + 302],mem_1_1[0 + 303],mem_1_1[0 + 304],mem_1_1[0 + 305],mem_1_1[0 + 306],mem_1_1[0 + 307],mem_1_1[0 + 308],mem_1_1[0 + 309],mem_1_1[0 + 310],mem_1_1[0 + 311],mem_1_1[0 + 312],mem_1_1[0 + 313],mem_1_1[0 + 314],mem_1_1[0 + 315],mem_1_1[0 + 316],mem_1_1[0 + 317],mem_1_1[0 + 318],mem_1_1[0 + 319],mem_1_1[0 + 320],mem_1_1[0 + 321],mem_1_1[0 + 322],mem_1_1[0 + 323],mem_1_1[0 + 324],mem_1_1[0 + 325],mem_1_1[0 + 326],mem_1_1[0 + 327],mem_1_1[0 + 328],mem_1_1[0 + 329],mem_1_1[0 + 330],mem_1_1[0 + 331],mem_1_1[0 + 332],mem_1_1[0 + 333],mem_1_1[0 + 334],mem_1_1[0 + 335],mem_1_1[0 + 336],mem_1_1[0 + 337],mem_1_1[0 + 338],mem_1_1[0 + 339],mem_1_1[0 + 340],mem_1_1[0 + 341],mem_1_1[0 + 342],mem_1_1[0 + 343],mem_1_1[0 + 344],mem_1_1[0 + 345],mem_1_1[0 + 346],mem_1_1[0 + 347],mem_1_1[0 + 348],mem_1_1[0 + 349],mem_1_1[0 + 350],mem_1_1[0 + 351],mem_1_1[0 + 352],mem_1_1[0 + 353],mem_1_1[0 + 354],mem_1_1[0 + 355],mem_1_1[0 + 356],mem_1_1[0 + 357],mem_1_1[0 + 358],mem_1_1[0 + 359],mem_1_1[0 + 360],mem_1_1[0 + 361],mem_1_1[0 + 362],mem_1_1[0 + 363],mem_1_1[0 + 364],mem_1_1[0 + 365],mem_1_1[0 + 366],mem_1_1[0 + 367],mem_1_1[0 + 368],mem_1_1[0 + 369],mem_1_1[0 + 370],mem_1_1[0 + 371],mem_1_1[0 + 372],mem_1_1[0 + 373],mem_1_1[0 + 374],mem_1_1[0 + 375],mem_1_1[0 + 376],mem_1_1[0 + 377],mem_1_1[0 + 378],mem_1_1[0 + 379],mem_1_1[0 + 380],mem_1_1[0 + 381],mem_1_1[0 + 382],mem_1_1[0 + 383],mem_1_1[0 + 384],mem_1_1[0 + 385],mem_1_1[0 + 386],mem_1_1[0 + 387],mem_1_1[0 + 388],mem_1_1[0 + 389],mem_1_1[0 + 390],mem_1_1[0 + 391],mem_1_1[0 + 392],mem_1_1[0 + 393],mem_1_1[0 + 394],mem_1_1[0 + 395],mem_1_1[0 + 396],mem_1_1[0 + 397],mem_1_1[0 + 398],mem_1_1[0 + 399],mem_1_1[0 + 400],mem_1_1[0 + 401],mem_1_1[0 + 402],mem_1_1[0 + 403],mem_1_1[0 + 404],mem_1_1[0 + 405],mem_1_1[0 + 406],mem_1_1[0 + 407],mem_1_1[0 + 408],mem_1_1[0 + 409],mem_1_1[0 + 410],mem_1_1[0 + 411],mem_1_1[0 + 412],mem_1_1[0 + 413],mem_1_1[0 + 414],mem_1_1[0 + 415],mem_1_1[0 + 416],mem_1_1[0 + 417],mem_1_1[0 + 418],mem_1_1[0 + 419],mem_1_1[0 + 420],mem_1_1[0 + 421],mem_1_1[0 + 422],mem_1_1[0 + 423],mem_1_1[0 + 424],mem_1_1[0 + 425],mem_1_1[0 + 426],mem_1_1[0 + 427],mem_1_1[0 + 428],mem_1_1[0 + 429],mem_1_1[0 + 430],mem_1_1[0 + 431],mem_1_1[0 + 432],mem_1_1[0 + 433],mem_1_1[0 + 434],mem_1_1[0 + 435],mem_1_1[0 + 436],mem_1_1[0 + 437],mem_1_1[0 + 438],mem_1_1[0 + 439],mem_1_1[0 + 440],mem_1_1[0 + 441],mem_1_1[0 + 442],mem_1_1[0 + 443],mem_1_1[0 + 444],mem_1_1[0 + 445],mem_1_1[0 + 446],mem_1_1[0 + 447],mem_1_1[0 + 448],mem_1_1[0 + 449],mem_1_1[0 + 450],mem_1_1[0 + 451],mem_1_1[0 + 452],mem_1_1[0 + 453],mem_1_1[0 + 454],mem_1_1[0 + 455],mem_1_1[0 + 456],mem_1_1[0 + 457],mem_1_1[0 + 458],mem_1_1[0 + 459],mem_1_1[0 + 460],mem_1_1[0 + 461],mem_1_1[0 + 462],mem_1_1[0 + 463],mem_1_1[0 + 464],mem_1_1[0 + 465],mem_1_1[0 + 466],mem_1_1[0 + 467],mem_1_1[0 + 468],mem_1_1[0 + 469],mem_1_1[0 + 470],mem_1_1[0 + 471],mem_1_1[0 + 472],mem_1_1[0 + 473],mem_1_1[0 + 474],mem_1_1[0 + 475],mem_1_1[0 + 476],mem_1_1[0 + 477],mem_1_1[0 + 478],mem_1_1[0 + 479],mem_1_1[0 + 480],mem_1_1[0 + 481],mem_1_1[0 + 482],mem_1_1[0 + 483],mem_1_1[0 + 484],mem_1_1[0 + 485],mem_1_1[0 + 486],mem_1_1[0 + 487],mem_1_1[0 + 488],mem_1_1[0 + 489],mem_1_1[0 + 490],mem_1_1[0 + 491],mem_1_1[0 + 492],mem_1_1[0 + 493],mem_1_1[0 + 494],mem_1_1[0 + 495],mem_1_1[0 + 496],mem_1_1[0 + 497],mem_1_1[0 + 498],mem_1_1[0 + 499],mem_1_1[0 + 500],mem_1_1[0 + 501],mem_1_1[0 + 502],mem_1_1[0 + 503],mem_1_1[0 + 504],mem_1_1[0 + 505],mem_1_1[0 + 506],mem_1_1[0 + 507],mem_1_1[0 + 508],mem_1_1[0 + 509],mem_1_1[0 + 510],mem_1_1[0 + 511],mem_1_1[0 + 512],mem_1_1[0 + 513],mem_1_1[0 + 514],mem_1_1[0 + 515],mem_1_1[0 + 516],mem_1_1[0 + 517],mem_1_1[0 + 518],mem_1_1[0 + 519],mem_1_1[0 + 520],mem_1_1[0 + 521],mem_1_1[0 + 522],mem_1_1[0 + 523],mem_1_1[0 + 524],mem_1_1[0 + 525],mem_1_1[0 + 526],mem_1_1[0 + 527],mem_1_1[0 + 528],mem_1_1[0 + 529],mem_1_1[0 + 530],mem_1_1[0 + 531],mem_1_1[0 + 532],mem_1_1[0 + 533],mem_1_1[0 + 534],mem_1_1[0 + 535],mem_1_1[0 + 536],mem_1_1[0 + 537],mem_1_1[0 + 538],mem_1_1[0 + 539],mem_1_1[0 + 540],mem_1_1[0 + 541],mem_1_1[0 + 542],mem_1_1[0 + 543],mem_1_1[0 + 544],mem_1_1[0 + 545],mem_1_1[0 + 546],mem_1_1[0 + 547],mem_1_1[0 + 548],mem_1_1[0 + 549],mem_1_1[0 + 550],mem_1_1[0 + 551],mem_1_1[0 + 552],mem_1_1[0 + 553],mem_1_1[0 + 554],mem_1_1[0 + 555],mem_1_1[0 + 556],mem_1_1[0 + 557],mem_1_1[0 + 558],mem_1_1[0 + 559],mem_1_1[0 + 560],mem_1_1[0 + 561],mem_1_1[0 + 562],mem_1_1[0 + 563],mem_1_1[0 + 564],mem_1_1[0 + 565],mem_1_1[0 + 566],mem_1_1[0 + 567],mem_1_1[0 + 568],mem_1_1[0 + 569],mem_1_1[0 + 570],mem_1_1[0 + 571],mem_1_1[0 + 572],mem_1_1[0 + 573],mem_1_1[0 + 574],mem_1_1[0 + 575],mem_1_1[0 + 576],mem_1_1[0 + 577],mem_1_1[0 + 578],mem_1_1[0 + 579],mem_1_1[0 + 580],mem_1_1[0 + 581],mem_1_1[0 + 582],mem_1_1[0 + 583],mem_1_1[0 + 584],mem_1_1[0 + 585],mem_1_1[0 + 586],mem_1_1[0 + 587],mem_1_1[0 + 588],mem_1_1[0 + 589],mem_1_1[0 + 590],mem_1_1[0 + 591],mem_1_1[0 + 592],mem_1_1[0 + 593],mem_1_1[0 + 594],mem_1_1[0 + 595],mem_1_1[0 + 596],mem_1_1[0 + 597],mem_1_1[0 + 598],mem_1_1[0 + 599],mem_1_1[0 + 600],mem_1_1[0 + 601],mem_1_1[0 + 602],mem_1_1[0 + 603],mem_1_1[0 + 604],mem_1_1[0 + 605],mem_1_1[0 + 606],mem_1_1[0 + 607],mem_1_1[0 + 608],mem_1_1[0 + 609],mem_1_1[0 + 610],mem_1_1[0 + 611],mem_1_1[0 + 612],mem_1_1[0 + 613],mem_1_1[0 + 614],mem_1_1[0 + 615],mem_1_1[0 + 616],mem_1_1[0 + 617],mem_1_1[0 + 618],mem_1_1[0 + 619],mem_1_1[0 + 620],mem_1_1[0 + 621],mem_1_1[0 + 622],mem_1_1[0 + 623],mem_1_1[0 + 624],mem_1_1[0 + 625],mem_1_1[0 + 626],mem_1_1[0 + 627],mem_1_1[0 + 628],mem_1_1[0 + 629],mem_1_1[0 + 630],mem_1_1[0 + 631],mem_1_1[0 + 632],mem_1_1[0 + 633],mem_1_1[0 + 634],mem_1_1[0 + 635],mem_1_1[0 + 636],mem_1_1[0 + 637],mem_1_1[0 + 638],mem_1_1[0 + 639],mem_1_1[0 + 640],mem_1_1[0 + 641],mem_1_1[0 + 642],mem_1_1[0 + 643],mem_1_1[0 + 644],mem_1_1[0 + 645],mem_1_1[0 + 646],mem_1_1[0 + 647],mem_1_1[0 + 648],mem_1_1[0 + 649],mem_1_1[0 + 650],mem_1_1[0 + 651],mem_1_1[0 + 652],mem_1_1[0 + 653],mem_1_1[0 + 654],mem_1_1[0 + 655],mem_1_1[0 + 656],mem_1_1[0 + 657],mem_1_1[0 + 658],mem_1_1[0 + 659],mem_1_1[0 + 660],mem_1_1[0 + 661],mem_1_1[0 + 662],mem_1_1[0 + 663],mem_1_1[0 + 664],mem_1_1[0 + 665],mem_1_1[0 + 666],mem_1_1[0 + 667],mem_1_1[0 + 668],mem_1_1[0 + 669],mem_1_1[0 + 670],mem_1_1[0 + 671],mem_1_1[0 + 672],mem_1_1[0 + 673],mem_1_1[0 + 674],mem_1_1[0 + 675],mem_1_1[0 + 676],mem_1_1[0 + 677],mem_1_1[0 + 678],mem_1_1[0 + 679],mem_1_1[0 + 680],mem_1_1[0 + 681],mem_1_1[0 + 682],mem_1_1[0 + 683],mem_1_1[0 + 684],mem_1_1[0 + 685],mem_1_1[0 + 686],mem_1_1[0 + 687],mem_1_1[0 + 688],mem_1_1[0 + 689],mem_1_1[0 + 690],mem_1_1[0 + 691],mem_1_1[0 + 692],mem_1_1[0 + 693],mem_1_1[0 + 694],mem_1_1[0 + 695],mem_1_1[0 + 696],mem_1_1[0 + 697],mem_1_1[0 + 698],mem_1_1[0 + 699],mem_1_1[0 + 700],mem_1_1[0 + 701],mem_1_1[0 + 702],mem_1_1[0 + 703],mem_1_1[0 + 704],mem_1_1[0 + 705],mem_1_1[0 + 706],mem_1_1[0 + 707],mem_1_1[0 + 708],mem_1_1[0 + 709],mem_1_1[0 + 710],mem_1_1[0 + 711],mem_1_1[0 + 712],mem_1_1[0 + 713],mem_1_1[0 + 714],mem_1_1[0 + 715],mem_1_1[0 + 716],mem_1_1[0 + 717],mem_1_1[0 + 718],mem_1_1[0 + 719],mem_1_1[0 + 720],mem_1_1[0 + 721],mem_1_1[0 + 722],mem_1_1[0 + 723],mem_1_1[0 + 724],mem_1_1[0 + 725],mem_1_1[0 + 726],mem_1_1[0 + 727],mem_1_1[0 + 728],mem_1_1[0 + 729],mem_1_1[0 + 730],mem_1_1[0 + 731],mem_1_1[0 + 732],mem_1_1[0 + 733],mem_1_1[0 + 734],mem_1_1[0 + 735],mem_1_1[0 + 736],mem_1_1[0 + 737],mem_1_1[0 + 738],mem_1_1[0 + 739],mem_1_1[0 + 740],mem_1_1[0 + 741],mem_1_1[0 + 742],mem_1_1[0 + 743],mem_1_1[0 + 744],mem_1_1[0 + 745],mem_1_1[0 + 746],mem_1_1[0 + 747],mem_1_1[0 + 748],mem_1_1[0 + 749],mem_1_1[0 + 750],mem_1_1[0 + 751],mem_1_1[0 + 752],mem_1_1[0 + 753],mem_1_1[0 + 754],mem_1_1[0 + 755],mem_1_1[0 + 756],mem_1_1[0 + 757],mem_1_1[0 + 758],mem_1_1[0 + 759],mem_1_1[0 + 760],mem_1_1[0 + 761],mem_1_1[0 + 762],mem_1_1[0 + 763],mem_1_1[0 + 764],mem_1_1[0 + 765],mem_1_1[0 + 766],mem_1_1[0 + 767],mem_1_1[0 + 768],mem_1_1[0 + 769],mem_1_1[0 + 770],mem_1_1[0 + 771],mem_1_1[0 + 772],mem_1_1[0 + 773],mem_1_1[0 + 774],mem_1_1[0 + 775],mem_1_1[0 + 776],mem_1_1[0 + 777],mem_1_1[0 + 778],mem_1_1[0 + 779],mem_1_1[0 + 780],mem_1_1[0 + 781],mem_1_1[0 + 782],mem_1_1[0 + 783],mem_1_1[0 + 784],mem_1_1[0 + 785],mem_1_1[0 + 786],mem_1_1[0 + 787],mem_1_1[0 + 788],mem_1_1[0 + 789],mem_1_1[0 + 790],mem_1_1[0 + 791],mem_1_1[0 + 792],mem_1_1[0 + 793],mem_1_1[0 + 794],mem_1_1[0 + 795],mem_1_1[0 + 796],mem_1_1[0 + 797],mem_1_1[0 + 798],mem_1_1[0 + 799],mem_1_1[0 + 800],mem_1_1[0 + 801],mem_1_1[0 + 802],mem_1_1[0 + 803],mem_1_1[0 + 804],mem_1_1[0 + 805],mem_1_1[0 + 806],mem_1_1[0 + 807],mem_1_1[0 + 808],mem_1_1[0 + 809],mem_1_1[0 + 810],mem_1_1[0 + 811],mem_1_1[0 + 812],mem_1_1[0 + 813],mem_1_1[0 + 814],mem_1_1[0 + 815],mem_1_1[0 + 816],mem_1_1[0 + 817],mem_1_1[0 + 818],mem_1_1[0 + 819],mem_1_1[0 + 820],mem_1_1[0 + 821],mem_1_1[0 + 822],mem_1_1[0 + 823],mem_1_1[0 + 824],mem_1_1[0 + 825],mem_1_1[0 + 826],mem_1_1[0 + 827],mem_1_1[0 + 828],mem_1_1[0 + 829],mem_1_1[0 + 830],mem_1_1[0 + 831],mem_1_1[0 + 832],mem_1_1[0 + 833],mem_1_1[0 + 834],mem_1_1[0 + 835],mem_1_1[0 + 836],mem_1_1[0 + 837],mem_1_1[0 + 838],mem_1_1[0 + 839],mem_1_1[0 + 840],mem_1_1[0 + 841],mem_1_1[0 + 842],mem_1_1[0 + 843],mem_1_1[0 + 844],mem_1_1[0 + 845],mem_1_1[0 + 846],mem_1_1[0 + 847],mem_1_1[0 + 848],mem_1_1[0 + 849],mem_1_1[0 + 850],mem_1_1[0 + 851],mem_1_1[0 + 852],mem_1_1[0 + 853],mem_1_1[0 + 854],mem_1_1[0 + 855],mem_1_1[0 + 856],mem_1_1[0 + 857],mem_1_1[0 + 858],mem_1_1[0 + 859],mem_1_1[0 + 860],mem_1_1[0 + 861],mem_1_1[0 + 862],mem_1_1[0 + 863],mem_1_1[0 + 864],mem_1_1[0 + 865],mem_1_1[0 + 866],mem_1_1[0 + 867],mem_1_1[0 + 868],mem_1_1[0 + 869],mem_1_1[0 + 870],mem_1_1[0 + 871],mem_1_1[0 + 872],mem_1_1[0 + 873],mem_1_1[0 + 874],mem_1_1[0 + 875],mem_1_1[0 + 876],mem_1_1[0 + 877],mem_1_1[0 + 878],mem_1_1[0 + 879],mem_1_1[0 + 880],mem_1_1[0 + 881],mem_1_1[0 + 882],mem_1_1[0 + 883],mem_1_1[0 + 884],mem_1_1[0 + 885],mem_1_1[0 + 886],mem_1_1[0 + 887],mem_1_1[0 + 888],mem_1_1[0 + 889],mem_1_1[0 + 890],mem_1_1[0 + 891],mem_1_1[0 + 892],mem_1_1[0 + 893],mem_1_1[0 + 894],mem_1_1[0 + 895],mem_1_1[0 + 896],mem_1_1[0 + 897],mem_1_1[0 + 898],mem_1_1[0 + 899],mem_1_1[0 + 900],mem_1_1[0 + 901],mem_1_1[0 + 902],mem_1_1[0 + 903],mem_1_1[0 + 904],mem_1_1[0 + 905],mem_1_1[0 + 906],mem_1_1[0 + 907],mem_1_1[0 + 908],mem_1_1[0 + 909],mem_1_1[0 + 910],mem_1_1[0 + 911],mem_1_1[0 + 912],mem_1_1[0 + 913],mem_1_1[0 + 914],mem_1_1[0 + 915],mem_1_1[0 + 916],mem_1_1[0 + 917],mem_1_1[0 + 918],mem_1_1[0 + 919],mem_1_1[0 + 920],mem_1_1[0 + 921],mem_1_1[0 + 922],mem_1_1[0 + 923],mem_1_1[0 + 924],mem_1_1[0 + 925],mem_1_1[0 + 926],mem_1_1[0 + 927],mem_1_1[0 + 928],mem_1_1[0 + 929],mem_1_1[0 + 930],mem_1_1[0 + 931],mem_1_1[0 + 932],mem_1_1[0 + 933],mem_1_1[0 + 934],mem_1_1[0 + 935],mem_1_1[0 + 936],mem_1_1[0 + 937],mem_1_1[0 + 938],mem_1_1[0 + 939],mem_1_1[0 + 940],mem_1_1[0 + 941],mem_1_1[0 + 942],mem_1_1[0 + 943],mem_1_1[0 + 944],mem_1_1[0 + 945],mem_1_1[0 + 946],mem_1_1[0 + 947],mem_1_1[0 + 948],mem_1_1[0 + 949],mem_1_1[0 + 950],mem_1_1[0 + 951],mem_1_1[0 + 952],mem_1_1[0 + 953],mem_1_1[0 + 954],mem_1_1[0 + 955],mem_1_1[0 + 956],mem_1_1[0 + 957],mem_1_1[0 + 958],mem_1_1[0 + 959],mem_1_1[0 + 960],mem_1_1[0 + 961],mem_1_1[0 + 962],mem_1_1[0 + 963],mem_1_1[0 + 964],mem_1_1[0 + 965],mem_1_1[0 + 966],mem_1_1[0 + 967],mem_1_1[0 + 968],mem_1_1[0 + 969],mem_1_1[0 + 970],mem_1_1[0 + 971],mem_1_1[0 + 972],mem_1_1[0 + 973],mem_1_1[0 + 974],mem_1_1[0 + 975],mem_1_1[0 + 976],mem_1_1[0 + 977],mem_1_1[0 + 978],mem_1_1[0 + 979],mem_1_1[0 + 980],mem_1_1[0 + 981],mem_1_1[0 + 982],mem_1_1[0 + 983],mem_1_1[0 + 984],mem_1_1[0 + 985],mem_1_1[0 + 986],mem_1_1[0 + 987],mem_1_1[0 + 988],mem_1_1[0 + 989],mem_1_1[0 + 990],mem_1_1[0 + 991],mem_1_1[0 + 992],mem_1_1[0 + 993],mem_1_1[0 + 994],mem_1_1[0 + 995],mem_1_1[0 + 996],mem_1_1[0 + 997],mem_1_1[0 + 998],mem_1_1[0 + 999],mem_1_1[0 + 1000],mem_1_1[0 + 1001],mem_1_1[0 + 1002],mem_1_1[0 + 1003],mem_1_1[0 + 1004],mem_1_1[0 + 1005],mem_1_1[0 + 1006],mem_1_1[0 + 1007],mem_1_1[0 + 1008],mem_1_1[0 + 1009],mem_1_1[0 + 1010],mem_1_1[0 + 1011],mem_1_1[0 + 1012],mem_1_1[0 + 1013],mem_1_1[0 + 1014],mem_1_1[0 + 1015],mem_1_1[0 + 1016],mem_1_1[0 + 1017],mem_1_1[0 + 1018],mem_1_1[0 + 1019],mem_1_1[0 + 1020],mem_1_1[0 + 1021],mem_1_1[0 + 1022],mem_1_1[0 + 1024 - 1] };
wire [8*(1024)-1:0] mem_2_1_flat_src;
assign mem_2_1_flat_src = {mem_2_1[0 + 0],mem_2_1[0 + 1],mem_2_1[0 + 2],mem_2_1[0 + 3],mem_2_1[0 + 4],mem_2_1[0 + 5],mem_2_1[0 + 6],mem_2_1[0 + 7],mem_2_1[0 + 8],mem_2_1[0 + 9],mem_2_1[0 + 10],mem_2_1[0 + 11],mem_2_1[0 + 12],mem_2_1[0 + 13],mem_2_1[0 + 14],mem_2_1[0 + 15],mem_2_1[0 + 16],mem_2_1[0 + 17],mem_2_1[0 + 18],mem_2_1[0 + 19],mem_2_1[0 + 20],mem_2_1[0 + 21],mem_2_1[0 + 22],mem_2_1[0 + 23],mem_2_1[0 + 24],mem_2_1[0 + 25],mem_2_1[0 + 26],mem_2_1[0 + 27],mem_2_1[0 + 28],mem_2_1[0 + 29],mem_2_1[0 + 30],mem_2_1[0 + 31],mem_2_1[0 + 32],mem_2_1[0 + 33],mem_2_1[0 + 34],mem_2_1[0 + 35],mem_2_1[0 + 36],mem_2_1[0 + 37],mem_2_1[0 + 38],mem_2_1[0 + 39],mem_2_1[0 + 40],mem_2_1[0 + 41],mem_2_1[0 + 42],mem_2_1[0 + 43],mem_2_1[0 + 44],mem_2_1[0 + 45],mem_2_1[0 + 46],mem_2_1[0 + 47],mem_2_1[0 + 48],mem_2_1[0 + 49],mem_2_1[0 + 50],mem_2_1[0 + 51],mem_2_1[0 + 52],mem_2_1[0 + 53],mem_2_1[0 + 54],mem_2_1[0 + 55],mem_2_1[0 + 56],mem_2_1[0 + 57],mem_2_1[0 + 58],mem_2_1[0 + 59],mem_2_1[0 + 60],mem_2_1[0 + 61],mem_2_1[0 + 62],mem_2_1[0 + 63],mem_2_1[0 + 64],mem_2_1[0 + 65],mem_2_1[0 + 66],mem_2_1[0 + 67],mem_2_1[0 + 68],mem_2_1[0 + 69],mem_2_1[0 + 70],mem_2_1[0 + 71],mem_2_1[0 + 72],mem_2_1[0 + 73],mem_2_1[0 + 74],mem_2_1[0 + 75],mem_2_1[0 + 76],mem_2_1[0 + 77],mem_2_1[0 + 78],mem_2_1[0 + 79],mem_2_1[0 + 80],mem_2_1[0 + 81],mem_2_1[0 + 82],mem_2_1[0 + 83],mem_2_1[0 + 84],mem_2_1[0 + 85],mem_2_1[0 + 86],mem_2_1[0 + 87],mem_2_1[0 + 88],mem_2_1[0 + 89],mem_2_1[0 + 90],mem_2_1[0 + 91],mem_2_1[0 + 92],mem_2_1[0 + 93],mem_2_1[0 + 94],mem_2_1[0 + 95],mem_2_1[0 + 96],mem_2_1[0 + 97],mem_2_1[0 + 98],mem_2_1[0 + 99],mem_2_1[0 + 100],mem_2_1[0 + 101],mem_2_1[0 + 102],mem_2_1[0 + 103],mem_2_1[0 + 104],mem_2_1[0 + 105],mem_2_1[0 + 106],mem_2_1[0 + 107],mem_2_1[0 + 108],mem_2_1[0 + 109],mem_2_1[0 + 110],mem_2_1[0 + 111],mem_2_1[0 + 112],mem_2_1[0 + 113],mem_2_1[0 + 114],mem_2_1[0 + 115],mem_2_1[0 + 116],mem_2_1[0 + 117],mem_2_1[0 + 118],mem_2_1[0 + 119],mem_2_1[0 + 120],mem_2_1[0 + 121],mem_2_1[0 + 122],mem_2_1[0 + 123],mem_2_1[0 + 124],mem_2_1[0 + 125],mem_2_1[0 + 126],mem_2_1[0 + 127],mem_2_1[0 + 128],mem_2_1[0 + 129],mem_2_1[0 + 130],mem_2_1[0 + 131],mem_2_1[0 + 132],mem_2_1[0 + 133],mem_2_1[0 + 134],mem_2_1[0 + 135],mem_2_1[0 + 136],mem_2_1[0 + 137],mem_2_1[0 + 138],mem_2_1[0 + 139],mem_2_1[0 + 140],mem_2_1[0 + 141],mem_2_1[0 + 142],mem_2_1[0 + 143],mem_2_1[0 + 144],mem_2_1[0 + 145],mem_2_1[0 + 146],mem_2_1[0 + 147],mem_2_1[0 + 148],mem_2_1[0 + 149],mem_2_1[0 + 150],mem_2_1[0 + 151],mem_2_1[0 + 152],mem_2_1[0 + 153],mem_2_1[0 + 154],mem_2_1[0 + 155],mem_2_1[0 + 156],mem_2_1[0 + 157],mem_2_1[0 + 158],mem_2_1[0 + 159],mem_2_1[0 + 160],mem_2_1[0 + 161],mem_2_1[0 + 162],mem_2_1[0 + 163],mem_2_1[0 + 164],mem_2_1[0 + 165],mem_2_1[0 + 166],mem_2_1[0 + 167],mem_2_1[0 + 168],mem_2_1[0 + 169],mem_2_1[0 + 170],mem_2_1[0 + 171],mem_2_1[0 + 172],mem_2_1[0 + 173],mem_2_1[0 + 174],mem_2_1[0 + 175],mem_2_1[0 + 176],mem_2_1[0 + 177],mem_2_1[0 + 178],mem_2_1[0 + 179],mem_2_1[0 + 180],mem_2_1[0 + 181],mem_2_1[0 + 182],mem_2_1[0 + 183],mem_2_1[0 + 184],mem_2_1[0 + 185],mem_2_1[0 + 186],mem_2_1[0 + 187],mem_2_1[0 + 188],mem_2_1[0 + 189],mem_2_1[0 + 190],mem_2_1[0 + 191],mem_2_1[0 + 192],mem_2_1[0 + 193],mem_2_1[0 + 194],mem_2_1[0 + 195],mem_2_1[0 + 196],mem_2_1[0 + 197],mem_2_1[0 + 198],mem_2_1[0 + 199],mem_2_1[0 + 200],mem_2_1[0 + 201],mem_2_1[0 + 202],mem_2_1[0 + 203],mem_2_1[0 + 204],mem_2_1[0 + 205],mem_2_1[0 + 206],mem_2_1[0 + 207],mem_2_1[0 + 208],mem_2_1[0 + 209],mem_2_1[0 + 210],mem_2_1[0 + 211],mem_2_1[0 + 212],mem_2_1[0 + 213],mem_2_1[0 + 214],mem_2_1[0 + 215],mem_2_1[0 + 216],mem_2_1[0 + 217],mem_2_1[0 + 218],mem_2_1[0 + 219],mem_2_1[0 + 220],mem_2_1[0 + 221],mem_2_1[0 + 222],mem_2_1[0 + 223],mem_2_1[0 + 224],mem_2_1[0 + 225],mem_2_1[0 + 226],mem_2_1[0 + 227],mem_2_1[0 + 228],mem_2_1[0 + 229],mem_2_1[0 + 230],mem_2_1[0 + 231],mem_2_1[0 + 232],mem_2_1[0 + 233],mem_2_1[0 + 234],mem_2_1[0 + 235],mem_2_1[0 + 236],mem_2_1[0 + 237],mem_2_1[0 + 238],mem_2_1[0 + 239],mem_2_1[0 + 240],mem_2_1[0 + 241],mem_2_1[0 + 242],mem_2_1[0 + 243],mem_2_1[0 + 244],mem_2_1[0 + 245],mem_2_1[0 + 246],mem_2_1[0 + 247],mem_2_1[0 + 248],mem_2_1[0 + 249],mem_2_1[0 + 250],mem_2_1[0 + 251],mem_2_1[0 + 252],mem_2_1[0 + 253],mem_2_1[0 + 254],mem_2_1[0 + 255],mem_2_1[0 + 256],mem_2_1[0 + 257],mem_2_1[0 + 258],mem_2_1[0 + 259],mem_2_1[0 + 260],mem_2_1[0 + 261],mem_2_1[0 + 262],mem_2_1[0 + 263],mem_2_1[0 + 264],mem_2_1[0 + 265],mem_2_1[0 + 266],mem_2_1[0 + 267],mem_2_1[0 + 268],mem_2_1[0 + 269],mem_2_1[0 + 270],mem_2_1[0 + 271],mem_2_1[0 + 272],mem_2_1[0 + 273],mem_2_1[0 + 274],mem_2_1[0 + 275],mem_2_1[0 + 276],mem_2_1[0 + 277],mem_2_1[0 + 278],mem_2_1[0 + 279],mem_2_1[0 + 280],mem_2_1[0 + 281],mem_2_1[0 + 282],mem_2_1[0 + 283],mem_2_1[0 + 284],mem_2_1[0 + 285],mem_2_1[0 + 286],mem_2_1[0 + 287],mem_2_1[0 + 288],mem_2_1[0 + 289],mem_2_1[0 + 290],mem_2_1[0 + 291],mem_2_1[0 + 292],mem_2_1[0 + 293],mem_2_1[0 + 294],mem_2_1[0 + 295],mem_2_1[0 + 296],mem_2_1[0 + 297],mem_2_1[0 + 298],mem_2_1[0 + 299],mem_2_1[0 + 300],mem_2_1[0 + 301],mem_2_1[0 + 302],mem_2_1[0 + 303],mem_2_1[0 + 304],mem_2_1[0 + 305],mem_2_1[0 + 306],mem_2_1[0 + 307],mem_2_1[0 + 308],mem_2_1[0 + 309],mem_2_1[0 + 310],mem_2_1[0 + 311],mem_2_1[0 + 312],mem_2_1[0 + 313],mem_2_1[0 + 314],mem_2_1[0 + 315],mem_2_1[0 + 316],mem_2_1[0 + 317],mem_2_1[0 + 318],mem_2_1[0 + 319],mem_2_1[0 + 320],mem_2_1[0 + 321],mem_2_1[0 + 322],mem_2_1[0 + 323],mem_2_1[0 + 324],mem_2_1[0 + 325],mem_2_1[0 + 326],mem_2_1[0 + 327],mem_2_1[0 + 328],mem_2_1[0 + 329],mem_2_1[0 + 330],mem_2_1[0 + 331],mem_2_1[0 + 332],mem_2_1[0 + 333],mem_2_1[0 + 334],mem_2_1[0 + 335],mem_2_1[0 + 336],mem_2_1[0 + 337],mem_2_1[0 + 338],mem_2_1[0 + 339],mem_2_1[0 + 340],mem_2_1[0 + 341],mem_2_1[0 + 342],mem_2_1[0 + 343],mem_2_1[0 + 344],mem_2_1[0 + 345],mem_2_1[0 + 346],mem_2_1[0 + 347],mem_2_1[0 + 348],mem_2_1[0 + 349],mem_2_1[0 + 350],mem_2_1[0 + 351],mem_2_1[0 + 352],mem_2_1[0 + 353],mem_2_1[0 + 354],mem_2_1[0 + 355],mem_2_1[0 + 356],mem_2_1[0 + 357],mem_2_1[0 + 358],mem_2_1[0 + 359],mem_2_1[0 + 360],mem_2_1[0 + 361],mem_2_1[0 + 362],mem_2_1[0 + 363],mem_2_1[0 + 364],mem_2_1[0 + 365],mem_2_1[0 + 366],mem_2_1[0 + 367],mem_2_1[0 + 368],mem_2_1[0 + 369],mem_2_1[0 + 370],mem_2_1[0 + 371],mem_2_1[0 + 372],mem_2_1[0 + 373],mem_2_1[0 + 374],mem_2_1[0 + 375],mem_2_1[0 + 376],mem_2_1[0 + 377],mem_2_1[0 + 378],mem_2_1[0 + 379],mem_2_1[0 + 380],mem_2_1[0 + 381],mem_2_1[0 + 382],mem_2_1[0 + 383],mem_2_1[0 + 384],mem_2_1[0 + 385],mem_2_1[0 + 386],mem_2_1[0 + 387],mem_2_1[0 + 388],mem_2_1[0 + 389],mem_2_1[0 + 390],mem_2_1[0 + 391],mem_2_1[0 + 392],mem_2_1[0 + 393],mem_2_1[0 + 394],mem_2_1[0 + 395],mem_2_1[0 + 396],mem_2_1[0 + 397],mem_2_1[0 + 398],mem_2_1[0 + 399],mem_2_1[0 + 400],mem_2_1[0 + 401],mem_2_1[0 + 402],mem_2_1[0 + 403],mem_2_1[0 + 404],mem_2_1[0 + 405],mem_2_1[0 + 406],mem_2_1[0 + 407],mem_2_1[0 + 408],mem_2_1[0 + 409],mem_2_1[0 + 410],mem_2_1[0 + 411],mem_2_1[0 + 412],mem_2_1[0 + 413],mem_2_1[0 + 414],mem_2_1[0 + 415],mem_2_1[0 + 416],mem_2_1[0 + 417],mem_2_1[0 + 418],mem_2_1[0 + 419],mem_2_1[0 + 420],mem_2_1[0 + 421],mem_2_1[0 + 422],mem_2_1[0 + 423],mem_2_1[0 + 424],mem_2_1[0 + 425],mem_2_1[0 + 426],mem_2_1[0 + 427],mem_2_1[0 + 428],mem_2_1[0 + 429],mem_2_1[0 + 430],mem_2_1[0 + 431],mem_2_1[0 + 432],mem_2_1[0 + 433],mem_2_1[0 + 434],mem_2_1[0 + 435],mem_2_1[0 + 436],mem_2_1[0 + 437],mem_2_1[0 + 438],mem_2_1[0 + 439],mem_2_1[0 + 440],mem_2_1[0 + 441],mem_2_1[0 + 442],mem_2_1[0 + 443],mem_2_1[0 + 444],mem_2_1[0 + 445],mem_2_1[0 + 446],mem_2_1[0 + 447],mem_2_1[0 + 448],mem_2_1[0 + 449],mem_2_1[0 + 450],mem_2_1[0 + 451],mem_2_1[0 + 452],mem_2_1[0 + 453],mem_2_1[0 + 454],mem_2_1[0 + 455],mem_2_1[0 + 456],mem_2_1[0 + 457],mem_2_1[0 + 458],mem_2_1[0 + 459],mem_2_1[0 + 460],mem_2_1[0 + 461],mem_2_1[0 + 462],mem_2_1[0 + 463],mem_2_1[0 + 464],mem_2_1[0 + 465],mem_2_1[0 + 466],mem_2_1[0 + 467],mem_2_1[0 + 468],mem_2_1[0 + 469],mem_2_1[0 + 470],mem_2_1[0 + 471],mem_2_1[0 + 472],mem_2_1[0 + 473],mem_2_1[0 + 474],mem_2_1[0 + 475],mem_2_1[0 + 476],mem_2_1[0 + 477],mem_2_1[0 + 478],mem_2_1[0 + 479],mem_2_1[0 + 480],mem_2_1[0 + 481],mem_2_1[0 + 482],mem_2_1[0 + 483],mem_2_1[0 + 484],mem_2_1[0 + 485],mem_2_1[0 + 486],mem_2_1[0 + 487],mem_2_1[0 + 488],mem_2_1[0 + 489],mem_2_1[0 + 490],mem_2_1[0 + 491],mem_2_1[0 + 492],mem_2_1[0 + 493],mem_2_1[0 + 494],mem_2_1[0 + 495],mem_2_1[0 + 496],mem_2_1[0 + 497],mem_2_1[0 + 498],mem_2_1[0 + 499],mem_2_1[0 + 500],mem_2_1[0 + 501],mem_2_1[0 + 502],mem_2_1[0 + 503],mem_2_1[0 + 504],mem_2_1[0 + 505],mem_2_1[0 + 506],mem_2_1[0 + 507],mem_2_1[0 + 508],mem_2_1[0 + 509],mem_2_1[0 + 510],mem_2_1[0 + 511],mem_2_1[0 + 512],mem_2_1[0 + 513],mem_2_1[0 + 514],mem_2_1[0 + 515],mem_2_1[0 + 516],mem_2_1[0 + 517],mem_2_1[0 + 518],mem_2_1[0 + 519],mem_2_1[0 + 520],mem_2_1[0 + 521],mem_2_1[0 + 522],mem_2_1[0 + 523],mem_2_1[0 + 524],mem_2_1[0 + 525],mem_2_1[0 + 526],mem_2_1[0 + 527],mem_2_1[0 + 528],mem_2_1[0 + 529],mem_2_1[0 + 530],mem_2_1[0 + 531],mem_2_1[0 + 532],mem_2_1[0 + 533],mem_2_1[0 + 534],mem_2_1[0 + 535],mem_2_1[0 + 536],mem_2_1[0 + 537],mem_2_1[0 + 538],mem_2_1[0 + 539],mem_2_1[0 + 540],mem_2_1[0 + 541],mem_2_1[0 + 542],mem_2_1[0 + 543],mem_2_1[0 + 544],mem_2_1[0 + 545],mem_2_1[0 + 546],mem_2_1[0 + 547],mem_2_1[0 + 548],mem_2_1[0 + 549],mem_2_1[0 + 550],mem_2_1[0 + 551],mem_2_1[0 + 552],mem_2_1[0 + 553],mem_2_1[0 + 554],mem_2_1[0 + 555],mem_2_1[0 + 556],mem_2_1[0 + 557],mem_2_1[0 + 558],mem_2_1[0 + 559],mem_2_1[0 + 560],mem_2_1[0 + 561],mem_2_1[0 + 562],mem_2_1[0 + 563],mem_2_1[0 + 564],mem_2_1[0 + 565],mem_2_1[0 + 566],mem_2_1[0 + 567],mem_2_1[0 + 568],mem_2_1[0 + 569],mem_2_1[0 + 570],mem_2_1[0 + 571],mem_2_1[0 + 572],mem_2_1[0 + 573],mem_2_1[0 + 574],mem_2_1[0 + 575],mem_2_1[0 + 576],mem_2_1[0 + 577],mem_2_1[0 + 578],mem_2_1[0 + 579],mem_2_1[0 + 580],mem_2_1[0 + 581],mem_2_1[0 + 582],mem_2_1[0 + 583],mem_2_1[0 + 584],mem_2_1[0 + 585],mem_2_1[0 + 586],mem_2_1[0 + 587],mem_2_1[0 + 588],mem_2_1[0 + 589],mem_2_1[0 + 590],mem_2_1[0 + 591],mem_2_1[0 + 592],mem_2_1[0 + 593],mem_2_1[0 + 594],mem_2_1[0 + 595],mem_2_1[0 + 596],mem_2_1[0 + 597],mem_2_1[0 + 598],mem_2_1[0 + 599],mem_2_1[0 + 600],mem_2_1[0 + 601],mem_2_1[0 + 602],mem_2_1[0 + 603],mem_2_1[0 + 604],mem_2_1[0 + 605],mem_2_1[0 + 606],mem_2_1[0 + 607],mem_2_1[0 + 608],mem_2_1[0 + 609],mem_2_1[0 + 610],mem_2_1[0 + 611],mem_2_1[0 + 612],mem_2_1[0 + 613],mem_2_1[0 + 614],mem_2_1[0 + 615],mem_2_1[0 + 616],mem_2_1[0 + 617],mem_2_1[0 + 618],mem_2_1[0 + 619],mem_2_1[0 + 620],mem_2_1[0 + 621],mem_2_1[0 + 622],mem_2_1[0 + 623],mem_2_1[0 + 624],mem_2_1[0 + 625],mem_2_1[0 + 626],mem_2_1[0 + 627],mem_2_1[0 + 628],mem_2_1[0 + 629],mem_2_1[0 + 630],mem_2_1[0 + 631],mem_2_1[0 + 632],mem_2_1[0 + 633],mem_2_1[0 + 634],mem_2_1[0 + 635],mem_2_1[0 + 636],mem_2_1[0 + 637],mem_2_1[0 + 638],mem_2_1[0 + 639],mem_2_1[0 + 640],mem_2_1[0 + 641],mem_2_1[0 + 642],mem_2_1[0 + 643],mem_2_1[0 + 644],mem_2_1[0 + 645],mem_2_1[0 + 646],mem_2_1[0 + 647],mem_2_1[0 + 648],mem_2_1[0 + 649],mem_2_1[0 + 650],mem_2_1[0 + 651],mem_2_1[0 + 652],mem_2_1[0 + 653],mem_2_1[0 + 654],mem_2_1[0 + 655],mem_2_1[0 + 656],mem_2_1[0 + 657],mem_2_1[0 + 658],mem_2_1[0 + 659],mem_2_1[0 + 660],mem_2_1[0 + 661],mem_2_1[0 + 662],mem_2_1[0 + 663],mem_2_1[0 + 664],mem_2_1[0 + 665],mem_2_1[0 + 666],mem_2_1[0 + 667],mem_2_1[0 + 668],mem_2_1[0 + 669],mem_2_1[0 + 670],mem_2_1[0 + 671],mem_2_1[0 + 672],mem_2_1[0 + 673],mem_2_1[0 + 674],mem_2_1[0 + 675],mem_2_1[0 + 676],mem_2_1[0 + 677],mem_2_1[0 + 678],mem_2_1[0 + 679],mem_2_1[0 + 680],mem_2_1[0 + 681],mem_2_1[0 + 682],mem_2_1[0 + 683],mem_2_1[0 + 684],mem_2_1[0 + 685],mem_2_1[0 + 686],mem_2_1[0 + 687],mem_2_1[0 + 688],mem_2_1[0 + 689],mem_2_1[0 + 690],mem_2_1[0 + 691],mem_2_1[0 + 692],mem_2_1[0 + 693],mem_2_1[0 + 694],mem_2_1[0 + 695],mem_2_1[0 + 696],mem_2_1[0 + 697],mem_2_1[0 + 698],mem_2_1[0 + 699],mem_2_1[0 + 700],mem_2_1[0 + 701],mem_2_1[0 + 702],mem_2_1[0 + 703],mem_2_1[0 + 704],mem_2_1[0 + 705],mem_2_1[0 + 706],mem_2_1[0 + 707],mem_2_1[0 + 708],mem_2_1[0 + 709],mem_2_1[0 + 710],mem_2_1[0 + 711],mem_2_1[0 + 712],mem_2_1[0 + 713],mem_2_1[0 + 714],mem_2_1[0 + 715],mem_2_1[0 + 716],mem_2_1[0 + 717],mem_2_1[0 + 718],mem_2_1[0 + 719],mem_2_1[0 + 720],mem_2_1[0 + 721],mem_2_1[0 + 722],mem_2_1[0 + 723],mem_2_1[0 + 724],mem_2_1[0 + 725],mem_2_1[0 + 726],mem_2_1[0 + 727],mem_2_1[0 + 728],mem_2_1[0 + 729],mem_2_1[0 + 730],mem_2_1[0 + 731],mem_2_1[0 + 732],mem_2_1[0 + 733],mem_2_1[0 + 734],mem_2_1[0 + 735],mem_2_1[0 + 736],mem_2_1[0 + 737],mem_2_1[0 + 738],mem_2_1[0 + 739],mem_2_1[0 + 740],mem_2_1[0 + 741],mem_2_1[0 + 742],mem_2_1[0 + 743],mem_2_1[0 + 744],mem_2_1[0 + 745],mem_2_1[0 + 746],mem_2_1[0 + 747],mem_2_1[0 + 748],mem_2_1[0 + 749],mem_2_1[0 + 750],mem_2_1[0 + 751],mem_2_1[0 + 752],mem_2_1[0 + 753],mem_2_1[0 + 754],mem_2_1[0 + 755],mem_2_1[0 + 756],mem_2_1[0 + 757],mem_2_1[0 + 758],mem_2_1[0 + 759],mem_2_1[0 + 760],mem_2_1[0 + 761],mem_2_1[0 + 762],mem_2_1[0 + 763],mem_2_1[0 + 764],mem_2_1[0 + 765],mem_2_1[0 + 766],mem_2_1[0 + 767],mem_2_1[0 + 768],mem_2_1[0 + 769],mem_2_1[0 + 770],mem_2_1[0 + 771],mem_2_1[0 + 772],mem_2_1[0 + 773],mem_2_1[0 + 774],mem_2_1[0 + 775],mem_2_1[0 + 776],mem_2_1[0 + 777],mem_2_1[0 + 778],mem_2_1[0 + 779],mem_2_1[0 + 780],mem_2_1[0 + 781],mem_2_1[0 + 782],mem_2_1[0 + 783],mem_2_1[0 + 784],mem_2_1[0 + 785],mem_2_1[0 + 786],mem_2_1[0 + 787],mem_2_1[0 + 788],mem_2_1[0 + 789],mem_2_1[0 + 790],mem_2_1[0 + 791],mem_2_1[0 + 792],mem_2_1[0 + 793],mem_2_1[0 + 794],mem_2_1[0 + 795],mem_2_1[0 + 796],mem_2_1[0 + 797],mem_2_1[0 + 798],mem_2_1[0 + 799],mem_2_1[0 + 800],mem_2_1[0 + 801],mem_2_1[0 + 802],mem_2_1[0 + 803],mem_2_1[0 + 804],mem_2_1[0 + 805],mem_2_1[0 + 806],mem_2_1[0 + 807],mem_2_1[0 + 808],mem_2_1[0 + 809],mem_2_1[0 + 810],mem_2_1[0 + 811],mem_2_1[0 + 812],mem_2_1[0 + 813],mem_2_1[0 + 814],mem_2_1[0 + 815],mem_2_1[0 + 816],mem_2_1[0 + 817],mem_2_1[0 + 818],mem_2_1[0 + 819],mem_2_1[0 + 820],mem_2_1[0 + 821],mem_2_1[0 + 822],mem_2_1[0 + 823],mem_2_1[0 + 824],mem_2_1[0 + 825],mem_2_1[0 + 826],mem_2_1[0 + 827],mem_2_1[0 + 828],mem_2_1[0 + 829],mem_2_1[0 + 830],mem_2_1[0 + 831],mem_2_1[0 + 832],mem_2_1[0 + 833],mem_2_1[0 + 834],mem_2_1[0 + 835],mem_2_1[0 + 836],mem_2_1[0 + 837],mem_2_1[0 + 838],mem_2_1[0 + 839],mem_2_1[0 + 840],mem_2_1[0 + 841],mem_2_1[0 + 842],mem_2_1[0 + 843],mem_2_1[0 + 844],mem_2_1[0 + 845],mem_2_1[0 + 846],mem_2_1[0 + 847],mem_2_1[0 + 848],mem_2_1[0 + 849],mem_2_1[0 + 850],mem_2_1[0 + 851],mem_2_1[0 + 852],mem_2_1[0 + 853],mem_2_1[0 + 854],mem_2_1[0 + 855],mem_2_1[0 + 856],mem_2_1[0 + 857],mem_2_1[0 + 858],mem_2_1[0 + 859],mem_2_1[0 + 860],mem_2_1[0 + 861],mem_2_1[0 + 862],mem_2_1[0 + 863],mem_2_1[0 + 864],mem_2_1[0 + 865],mem_2_1[0 + 866],mem_2_1[0 + 867],mem_2_1[0 + 868],mem_2_1[0 + 869],mem_2_1[0 + 870],mem_2_1[0 + 871],mem_2_1[0 + 872],mem_2_1[0 + 873],mem_2_1[0 + 874],mem_2_1[0 + 875],mem_2_1[0 + 876],mem_2_1[0 + 877],mem_2_1[0 + 878],mem_2_1[0 + 879],mem_2_1[0 + 880],mem_2_1[0 + 881],mem_2_1[0 + 882],mem_2_1[0 + 883],mem_2_1[0 + 884],mem_2_1[0 + 885],mem_2_1[0 + 886],mem_2_1[0 + 887],mem_2_1[0 + 888],mem_2_1[0 + 889],mem_2_1[0 + 890],mem_2_1[0 + 891],mem_2_1[0 + 892],mem_2_1[0 + 893],mem_2_1[0 + 894],mem_2_1[0 + 895],mem_2_1[0 + 896],mem_2_1[0 + 897],mem_2_1[0 + 898],mem_2_1[0 + 899],mem_2_1[0 + 900],mem_2_1[0 + 901],mem_2_1[0 + 902],mem_2_1[0 + 903],mem_2_1[0 + 904],mem_2_1[0 + 905],mem_2_1[0 + 906],mem_2_1[0 + 907],mem_2_1[0 + 908],mem_2_1[0 + 909],mem_2_1[0 + 910],mem_2_1[0 + 911],mem_2_1[0 + 912],mem_2_1[0 + 913],mem_2_1[0 + 914],mem_2_1[0 + 915],mem_2_1[0 + 916],mem_2_1[0 + 917],mem_2_1[0 + 918],mem_2_1[0 + 919],mem_2_1[0 + 920],mem_2_1[0 + 921],mem_2_1[0 + 922],mem_2_1[0 + 923],mem_2_1[0 + 924],mem_2_1[0 + 925],mem_2_1[0 + 926],mem_2_1[0 + 927],mem_2_1[0 + 928],mem_2_1[0 + 929],mem_2_1[0 + 930],mem_2_1[0 + 931],mem_2_1[0 + 932],mem_2_1[0 + 933],mem_2_1[0 + 934],mem_2_1[0 + 935],mem_2_1[0 + 936],mem_2_1[0 + 937],mem_2_1[0 + 938],mem_2_1[0 + 939],mem_2_1[0 + 940],mem_2_1[0 + 941],mem_2_1[0 + 942],mem_2_1[0 + 943],mem_2_1[0 + 944],mem_2_1[0 + 945],mem_2_1[0 + 946],mem_2_1[0 + 947],mem_2_1[0 + 948],mem_2_1[0 + 949],mem_2_1[0 + 950],mem_2_1[0 + 951],mem_2_1[0 + 952],mem_2_1[0 + 953],mem_2_1[0 + 954],mem_2_1[0 + 955],mem_2_1[0 + 956],mem_2_1[0 + 957],mem_2_1[0 + 958],mem_2_1[0 + 959],mem_2_1[0 + 960],mem_2_1[0 + 961],mem_2_1[0 + 962],mem_2_1[0 + 963],mem_2_1[0 + 964],mem_2_1[0 + 965],mem_2_1[0 + 966],mem_2_1[0 + 967],mem_2_1[0 + 968],mem_2_1[0 + 969],mem_2_1[0 + 970],mem_2_1[0 + 971],mem_2_1[0 + 972],mem_2_1[0 + 973],mem_2_1[0 + 974],mem_2_1[0 + 975],mem_2_1[0 + 976],mem_2_1[0 + 977],mem_2_1[0 + 978],mem_2_1[0 + 979],mem_2_1[0 + 980],mem_2_1[0 + 981],mem_2_1[0 + 982],mem_2_1[0 + 983],mem_2_1[0 + 984],mem_2_1[0 + 985],mem_2_1[0 + 986],mem_2_1[0 + 987],mem_2_1[0 + 988],mem_2_1[0 + 989],mem_2_1[0 + 990],mem_2_1[0 + 991],mem_2_1[0 + 992],mem_2_1[0 + 993],mem_2_1[0 + 994],mem_2_1[0 + 995],mem_2_1[0 + 996],mem_2_1[0 + 997],mem_2_1[0 + 998],mem_2_1[0 + 999],mem_2_1[0 + 1000],mem_2_1[0 + 1001],mem_2_1[0 + 1002],mem_2_1[0 + 1003],mem_2_1[0 + 1004],mem_2_1[0 + 1005],mem_2_1[0 + 1006],mem_2_1[0 + 1007],mem_2_1[0 + 1008],mem_2_1[0 + 1009],mem_2_1[0 + 1010],mem_2_1[0 + 1011],mem_2_1[0 + 1012],mem_2_1[0 + 1013],mem_2_1[0 + 1014],mem_2_1[0 + 1015],mem_2_1[0 + 1016],mem_2_1[0 + 1017],mem_2_1[0 + 1018],mem_2_1[0 + 1019],mem_2_1[0 + 1020],mem_2_1[0 + 1021],mem_2_1[0 + 1022],mem_2_1[0 + 1024 - 1] };
wire [8*(1024)-1:0] mem_3_1_flat_src;
assign mem_3_1_flat_src = {mem_3_1[0 + 0],mem_3_1[0 + 1],mem_3_1[0 + 2],mem_3_1[0 + 3],mem_3_1[0 + 4],mem_3_1[0 + 5],mem_3_1[0 + 6],mem_3_1[0 + 7],mem_3_1[0 + 8],mem_3_1[0 + 9],mem_3_1[0 + 10],mem_3_1[0 + 11],mem_3_1[0 + 12],mem_3_1[0 + 13],mem_3_1[0 + 14],mem_3_1[0 + 15],mem_3_1[0 + 16],mem_3_1[0 + 17],mem_3_1[0 + 18],mem_3_1[0 + 19],mem_3_1[0 + 20],mem_3_1[0 + 21],mem_3_1[0 + 22],mem_3_1[0 + 23],mem_3_1[0 + 24],mem_3_1[0 + 25],mem_3_1[0 + 26],mem_3_1[0 + 27],mem_3_1[0 + 28],mem_3_1[0 + 29],mem_3_1[0 + 30],mem_3_1[0 + 31],mem_3_1[0 + 32],mem_3_1[0 + 33],mem_3_1[0 + 34],mem_3_1[0 + 35],mem_3_1[0 + 36],mem_3_1[0 + 37],mem_3_1[0 + 38],mem_3_1[0 + 39],mem_3_1[0 + 40],mem_3_1[0 + 41],mem_3_1[0 + 42],mem_3_1[0 + 43],mem_3_1[0 + 44],mem_3_1[0 + 45],mem_3_1[0 + 46],mem_3_1[0 + 47],mem_3_1[0 + 48],mem_3_1[0 + 49],mem_3_1[0 + 50],mem_3_1[0 + 51],mem_3_1[0 + 52],mem_3_1[0 + 53],mem_3_1[0 + 54],mem_3_1[0 + 55],mem_3_1[0 + 56],mem_3_1[0 + 57],mem_3_1[0 + 58],mem_3_1[0 + 59],mem_3_1[0 + 60],mem_3_1[0 + 61],mem_3_1[0 + 62],mem_3_1[0 + 63],mem_3_1[0 + 64],mem_3_1[0 + 65],mem_3_1[0 + 66],mem_3_1[0 + 67],mem_3_1[0 + 68],mem_3_1[0 + 69],mem_3_1[0 + 70],mem_3_1[0 + 71],mem_3_1[0 + 72],mem_3_1[0 + 73],mem_3_1[0 + 74],mem_3_1[0 + 75],mem_3_1[0 + 76],mem_3_1[0 + 77],mem_3_1[0 + 78],mem_3_1[0 + 79],mem_3_1[0 + 80],mem_3_1[0 + 81],mem_3_1[0 + 82],mem_3_1[0 + 83],mem_3_1[0 + 84],mem_3_1[0 + 85],mem_3_1[0 + 86],mem_3_1[0 + 87],mem_3_1[0 + 88],mem_3_1[0 + 89],mem_3_1[0 + 90],mem_3_1[0 + 91],mem_3_1[0 + 92],mem_3_1[0 + 93],mem_3_1[0 + 94],mem_3_1[0 + 95],mem_3_1[0 + 96],mem_3_1[0 + 97],mem_3_1[0 + 98],mem_3_1[0 + 99],mem_3_1[0 + 100],mem_3_1[0 + 101],mem_3_1[0 + 102],mem_3_1[0 + 103],mem_3_1[0 + 104],mem_3_1[0 + 105],mem_3_1[0 + 106],mem_3_1[0 + 107],mem_3_1[0 + 108],mem_3_1[0 + 109],mem_3_1[0 + 110],mem_3_1[0 + 111],mem_3_1[0 + 112],mem_3_1[0 + 113],mem_3_1[0 + 114],mem_3_1[0 + 115],mem_3_1[0 + 116],mem_3_1[0 + 117],mem_3_1[0 + 118],mem_3_1[0 + 119],mem_3_1[0 + 120],mem_3_1[0 + 121],mem_3_1[0 + 122],mem_3_1[0 + 123],mem_3_1[0 + 124],mem_3_1[0 + 125],mem_3_1[0 + 126],mem_3_1[0 + 127],mem_3_1[0 + 128],mem_3_1[0 + 129],mem_3_1[0 + 130],mem_3_1[0 + 131],mem_3_1[0 + 132],mem_3_1[0 + 133],mem_3_1[0 + 134],mem_3_1[0 + 135],mem_3_1[0 + 136],mem_3_1[0 + 137],mem_3_1[0 + 138],mem_3_1[0 + 139],mem_3_1[0 + 140],mem_3_1[0 + 141],mem_3_1[0 + 142],mem_3_1[0 + 143],mem_3_1[0 + 144],mem_3_1[0 + 145],mem_3_1[0 + 146],mem_3_1[0 + 147],mem_3_1[0 + 148],mem_3_1[0 + 149],mem_3_1[0 + 150],mem_3_1[0 + 151],mem_3_1[0 + 152],mem_3_1[0 + 153],mem_3_1[0 + 154],mem_3_1[0 + 155],mem_3_1[0 + 156],mem_3_1[0 + 157],mem_3_1[0 + 158],mem_3_1[0 + 159],mem_3_1[0 + 160],mem_3_1[0 + 161],mem_3_1[0 + 162],mem_3_1[0 + 163],mem_3_1[0 + 164],mem_3_1[0 + 165],mem_3_1[0 + 166],mem_3_1[0 + 167],mem_3_1[0 + 168],mem_3_1[0 + 169],mem_3_1[0 + 170],mem_3_1[0 + 171],mem_3_1[0 + 172],mem_3_1[0 + 173],mem_3_1[0 + 174],mem_3_1[0 + 175],mem_3_1[0 + 176],mem_3_1[0 + 177],mem_3_1[0 + 178],mem_3_1[0 + 179],mem_3_1[0 + 180],mem_3_1[0 + 181],mem_3_1[0 + 182],mem_3_1[0 + 183],mem_3_1[0 + 184],mem_3_1[0 + 185],mem_3_1[0 + 186],mem_3_1[0 + 187],mem_3_1[0 + 188],mem_3_1[0 + 189],mem_3_1[0 + 190],mem_3_1[0 + 191],mem_3_1[0 + 192],mem_3_1[0 + 193],mem_3_1[0 + 194],mem_3_1[0 + 195],mem_3_1[0 + 196],mem_3_1[0 + 197],mem_3_1[0 + 198],mem_3_1[0 + 199],mem_3_1[0 + 200],mem_3_1[0 + 201],mem_3_1[0 + 202],mem_3_1[0 + 203],mem_3_1[0 + 204],mem_3_1[0 + 205],mem_3_1[0 + 206],mem_3_1[0 + 207],mem_3_1[0 + 208],mem_3_1[0 + 209],mem_3_1[0 + 210],mem_3_1[0 + 211],mem_3_1[0 + 212],mem_3_1[0 + 213],mem_3_1[0 + 214],mem_3_1[0 + 215],mem_3_1[0 + 216],mem_3_1[0 + 217],mem_3_1[0 + 218],mem_3_1[0 + 219],mem_3_1[0 + 220],mem_3_1[0 + 221],mem_3_1[0 + 222],mem_3_1[0 + 223],mem_3_1[0 + 224],mem_3_1[0 + 225],mem_3_1[0 + 226],mem_3_1[0 + 227],mem_3_1[0 + 228],mem_3_1[0 + 229],mem_3_1[0 + 230],mem_3_1[0 + 231],mem_3_1[0 + 232],mem_3_1[0 + 233],mem_3_1[0 + 234],mem_3_1[0 + 235],mem_3_1[0 + 236],mem_3_1[0 + 237],mem_3_1[0 + 238],mem_3_1[0 + 239],mem_3_1[0 + 240],mem_3_1[0 + 241],mem_3_1[0 + 242],mem_3_1[0 + 243],mem_3_1[0 + 244],mem_3_1[0 + 245],mem_3_1[0 + 246],mem_3_1[0 + 247],mem_3_1[0 + 248],mem_3_1[0 + 249],mem_3_1[0 + 250],mem_3_1[0 + 251],mem_3_1[0 + 252],mem_3_1[0 + 253],mem_3_1[0 + 254],mem_3_1[0 + 255],mem_3_1[0 + 256],mem_3_1[0 + 257],mem_3_1[0 + 258],mem_3_1[0 + 259],mem_3_1[0 + 260],mem_3_1[0 + 261],mem_3_1[0 + 262],mem_3_1[0 + 263],mem_3_1[0 + 264],mem_3_1[0 + 265],mem_3_1[0 + 266],mem_3_1[0 + 267],mem_3_1[0 + 268],mem_3_1[0 + 269],mem_3_1[0 + 270],mem_3_1[0 + 271],mem_3_1[0 + 272],mem_3_1[0 + 273],mem_3_1[0 + 274],mem_3_1[0 + 275],mem_3_1[0 + 276],mem_3_1[0 + 277],mem_3_1[0 + 278],mem_3_1[0 + 279],mem_3_1[0 + 280],mem_3_1[0 + 281],mem_3_1[0 + 282],mem_3_1[0 + 283],mem_3_1[0 + 284],mem_3_1[0 + 285],mem_3_1[0 + 286],mem_3_1[0 + 287],mem_3_1[0 + 288],mem_3_1[0 + 289],mem_3_1[0 + 290],mem_3_1[0 + 291],mem_3_1[0 + 292],mem_3_1[0 + 293],mem_3_1[0 + 294],mem_3_1[0 + 295],mem_3_1[0 + 296],mem_3_1[0 + 297],mem_3_1[0 + 298],mem_3_1[0 + 299],mem_3_1[0 + 300],mem_3_1[0 + 301],mem_3_1[0 + 302],mem_3_1[0 + 303],mem_3_1[0 + 304],mem_3_1[0 + 305],mem_3_1[0 + 306],mem_3_1[0 + 307],mem_3_1[0 + 308],mem_3_1[0 + 309],mem_3_1[0 + 310],mem_3_1[0 + 311],mem_3_1[0 + 312],mem_3_1[0 + 313],mem_3_1[0 + 314],mem_3_1[0 + 315],mem_3_1[0 + 316],mem_3_1[0 + 317],mem_3_1[0 + 318],mem_3_1[0 + 319],mem_3_1[0 + 320],mem_3_1[0 + 321],mem_3_1[0 + 322],mem_3_1[0 + 323],mem_3_1[0 + 324],mem_3_1[0 + 325],mem_3_1[0 + 326],mem_3_1[0 + 327],mem_3_1[0 + 328],mem_3_1[0 + 329],mem_3_1[0 + 330],mem_3_1[0 + 331],mem_3_1[0 + 332],mem_3_1[0 + 333],mem_3_1[0 + 334],mem_3_1[0 + 335],mem_3_1[0 + 336],mem_3_1[0 + 337],mem_3_1[0 + 338],mem_3_1[0 + 339],mem_3_1[0 + 340],mem_3_1[0 + 341],mem_3_1[0 + 342],mem_3_1[0 + 343],mem_3_1[0 + 344],mem_3_1[0 + 345],mem_3_1[0 + 346],mem_3_1[0 + 347],mem_3_1[0 + 348],mem_3_1[0 + 349],mem_3_1[0 + 350],mem_3_1[0 + 351],mem_3_1[0 + 352],mem_3_1[0 + 353],mem_3_1[0 + 354],mem_3_1[0 + 355],mem_3_1[0 + 356],mem_3_1[0 + 357],mem_3_1[0 + 358],mem_3_1[0 + 359],mem_3_1[0 + 360],mem_3_1[0 + 361],mem_3_1[0 + 362],mem_3_1[0 + 363],mem_3_1[0 + 364],mem_3_1[0 + 365],mem_3_1[0 + 366],mem_3_1[0 + 367],mem_3_1[0 + 368],mem_3_1[0 + 369],mem_3_1[0 + 370],mem_3_1[0 + 371],mem_3_1[0 + 372],mem_3_1[0 + 373],mem_3_1[0 + 374],mem_3_1[0 + 375],mem_3_1[0 + 376],mem_3_1[0 + 377],mem_3_1[0 + 378],mem_3_1[0 + 379],mem_3_1[0 + 380],mem_3_1[0 + 381],mem_3_1[0 + 382],mem_3_1[0 + 383],mem_3_1[0 + 384],mem_3_1[0 + 385],mem_3_1[0 + 386],mem_3_1[0 + 387],mem_3_1[0 + 388],mem_3_1[0 + 389],mem_3_1[0 + 390],mem_3_1[0 + 391],mem_3_1[0 + 392],mem_3_1[0 + 393],mem_3_1[0 + 394],mem_3_1[0 + 395],mem_3_1[0 + 396],mem_3_1[0 + 397],mem_3_1[0 + 398],mem_3_1[0 + 399],mem_3_1[0 + 400],mem_3_1[0 + 401],mem_3_1[0 + 402],mem_3_1[0 + 403],mem_3_1[0 + 404],mem_3_1[0 + 405],mem_3_1[0 + 406],mem_3_1[0 + 407],mem_3_1[0 + 408],mem_3_1[0 + 409],mem_3_1[0 + 410],mem_3_1[0 + 411],mem_3_1[0 + 412],mem_3_1[0 + 413],mem_3_1[0 + 414],mem_3_1[0 + 415],mem_3_1[0 + 416],mem_3_1[0 + 417],mem_3_1[0 + 418],mem_3_1[0 + 419],mem_3_1[0 + 420],mem_3_1[0 + 421],mem_3_1[0 + 422],mem_3_1[0 + 423],mem_3_1[0 + 424],mem_3_1[0 + 425],mem_3_1[0 + 426],mem_3_1[0 + 427],mem_3_1[0 + 428],mem_3_1[0 + 429],mem_3_1[0 + 430],mem_3_1[0 + 431],mem_3_1[0 + 432],mem_3_1[0 + 433],mem_3_1[0 + 434],mem_3_1[0 + 435],mem_3_1[0 + 436],mem_3_1[0 + 437],mem_3_1[0 + 438],mem_3_1[0 + 439],mem_3_1[0 + 440],mem_3_1[0 + 441],mem_3_1[0 + 442],mem_3_1[0 + 443],mem_3_1[0 + 444],mem_3_1[0 + 445],mem_3_1[0 + 446],mem_3_1[0 + 447],mem_3_1[0 + 448],mem_3_1[0 + 449],mem_3_1[0 + 450],mem_3_1[0 + 451],mem_3_1[0 + 452],mem_3_1[0 + 453],mem_3_1[0 + 454],mem_3_1[0 + 455],mem_3_1[0 + 456],mem_3_1[0 + 457],mem_3_1[0 + 458],mem_3_1[0 + 459],mem_3_1[0 + 460],mem_3_1[0 + 461],mem_3_1[0 + 462],mem_3_1[0 + 463],mem_3_1[0 + 464],mem_3_1[0 + 465],mem_3_1[0 + 466],mem_3_1[0 + 467],mem_3_1[0 + 468],mem_3_1[0 + 469],mem_3_1[0 + 470],mem_3_1[0 + 471],mem_3_1[0 + 472],mem_3_1[0 + 473],mem_3_1[0 + 474],mem_3_1[0 + 475],mem_3_1[0 + 476],mem_3_1[0 + 477],mem_3_1[0 + 478],mem_3_1[0 + 479],mem_3_1[0 + 480],mem_3_1[0 + 481],mem_3_1[0 + 482],mem_3_1[0 + 483],mem_3_1[0 + 484],mem_3_1[0 + 485],mem_3_1[0 + 486],mem_3_1[0 + 487],mem_3_1[0 + 488],mem_3_1[0 + 489],mem_3_1[0 + 490],mem_3_1[0 + 491],mem_3_1[0 + 492],mem_3_1[0 + 493],mem_3_1[0 + 494],mem_3_1[0 + 495],mem_3_1[0 + 496],mem_3_1[0 + 497],mem_3_1[0 + 498],mem_3_1[0 + 499],mem_3_1[0 + 500],mem_3_1[0 + 501],mem_3_1[0 + 502],mem_3_1[0 + 503],mem_3_1[0 + 504],mem_3_1[0 + 505],mem_3_1[0 + 506],mem_3_1[0 + 507],mem_3_1[0 + 508],mem_3_1[0 + 509],mem_3_1[0 + 510],mem_3_1[0 + 511],mem_3_1[0 + 512],mem_3_1[0 + 513],mem_3_1[0 + 514],mem_3_1[0 + 515],mem_3_1[0 + 516],mem_3_1[0 + 517],mem_3_1[0 + 518],mem_3_1[0 + 519],mem_3_1[0 + 520],mem_3_1[0 + 521],mem_3_1[0 + 522],mem_3_1[0 + 523],mem_3_1[0 + 524],mem_3_1[0 + 525],mem_3_1[0 + 526],mem_3_1[0 + 527],mem_3_1[0 + 528],mem_3_1[0 + 529],mem_3_1[0 + 530],mem_3_1[0 + 531],mem_3_1[0 + 532],mem_3_1[0 + 533],mem_3_1[0 + 534],mem_3_1[0 + 535],mem_3_1[0 + 536],mem_3_1[0 + 537],mem_3_1[0 + 538],mem_3_1[0 + 539],mem_3_1[0 + 540],mem_3_1[0 + 541],mem_3_1[0 + 542],mem_3_1[0 + 543],mem_3_1[0 + 544],mem_3_1[0 + 545],mem_3_1[0 + 546],mem_3_1[0 + 547],mem_3_1[0 + 548],mem_3_1[0 + 549],mem_3_1[0 + 550],mem_3_1[0 + 551],mem_3_1[0 + 552],mem_3_1[0 + 553],mem_3_1[0 + 554],mem_3_1[0 + 555],mem_3_1[0 + 556],mem_3_1[0 + 557],mem_3_1[0 + 558],mem_3_1[0 + 559],mem_3_1[0 + 560],mem_3_1[0 + 561],mem_3_1[0 + 562],mem_3_1[0 + 563],mem_3_1[0 + 564],mem_3_1[0 + 565],mem_3_1[0 + 566],mem_3_1[0 + 567],mem_3_1[0 + 568],mem_3_1[0 + 569],mem_3_1[0 + 570],mem_3_1[0 + 571],mem_3_1[0 + 572],mem_3_1[0 + 573],mem_3_1[0 + 574],mem_3_1[0 + 575],mem_3_1[0 + 576],mem_3_1[0 + 577],mem_3_1[0 + 578],mem_3_1[0 + 579],mem_3_1[0 + 580],mem_3_1[0 + 581],mem_3_1[0 + 582],mem_3_1[0 + 583],mem_3_1[0 + 584],mem_3_1[0 + 585],mem_3_1[0 + 586],mem_3_1[0 + 587],mem_3_1[0 + 588],mem_3_1[0 + 589],mem_3_1[0 + 590],mem_3_1[0 + 591],mem_3_1[0 + 592],mem_3_1[0 + 593],mem_3_1[0 + 594],mem_3_1[0 + 595],mem_3_1[0 + 596],mem_3_1[0 + 597],mem_3_1[0 + 598],mem_3_1[0 + 599],mem_3_1[0 + 600],mem_3_1[0 + 601],mem_3_1[0 + 602],mem_3_1[0 + 603],mem_3_1[0 + 604],mem_3_1[0 + 605],mem_3_1[0 + 606],mem_3_1[0 + 607],mem_3_1[0 + 608],mem_3_1[0 + 609],mem_3_1[0 + 610],mem_3_1[0 + 611],mem_3_1[0 + 612],mem_3_1[0 + 613],mem_3_1[0 + 614],mem_3_1[0 + 615],mem_3_1[0 + 616],mem_3_1[0 + 617],mem_3_1[0 + 618],mem_3_1[0 + 619],mem_3_1[0 + 620],mem_3_1[0 + 621],mem_3_1[0 + 622],mem_3_1[0 + 623],mem_3_1[0 + 624],mem_3_1[0 + 625],mem_3_1[0 + 626],mem_3_1[0 + 627],mem_3_1[0 + 628],mem_3_1[0 + 629],mem_3_1[0 + 630],mem_3_1[0 + 631],mem_3_1[0 + 632],mem_3_1[0 + 633],mem_3_1[0 + 634],mem_3_1[0 + 635],mem_3_1[0 + 636],mem_3_1[0 + 637],mem_3_1[0 + 638],mem_3_1[0 + 639],mem_3_1[0 + 640],mem_3_1[0 + 641],mem_3_1[0 + 642],mem_3_1[0 + 643],mem_3_1[0 + 644],mem_3_1[0 + 645],mem_3_1[0 + 646],mem_3_1[0 + 647],mem_3_1[0 + 648],mem_3_1[0 + 649],mem_3_1[0 + 650],mem_3_1[0 + 651],mem_3_1[0 + 652],mem_3_1[0 + 653],mem_3_1[0 + 654],mem_3_1[0 + 655],mem_3_1[0 + 656],mem_3_1[0 + 657],mem_3_1[0 + 658],mem_3_1[0 + 659],mem_3_1[0 + 660],mem_3_1[0 + 661],mem_3_1[0 + 662],mem_3_1[0 + 663],mem_3_1[0 + 664],mem_3_1[0 + 665],mem_3_1[0 + 666],mem_3_1[0 + 667],mem_3_1[0 + 668],mem_3_1[0 + 669],mem_3_1[0 + 670],mem_3_1[0 + 671],mem_3_1[0 + 672],mem_3_1[0 + 673],mem_3_1[0 + 674],mem_3_1[0 + 675],mem_3_1[0 + 676],mem_3_1[0 + 677],mem_3_1[0 + 678],mem_3_1[0 + 679],mem_3_1[0 + 680],mem_3_1[0 + 681],mem_3_1[0 + 682],mem_3_1[0 + 683],mem_3_1[0 + 684],mem_3_1[0 + 685],mem_3_1[0 + 686],mem_3_1[0 + 687],mem_3_1[0 + 688],mem_3_1[0 + 689],mem_3_1[0 + 690],mem_3_1[0 + 691],mem_3_1[0 + 692],mem_3_1[0 + 693],mem_3_1[0 + 694],mem_3_1[0 + 695],mem_3_1[0 + 696],mem_3_1[0 + 697],mem_3_1[0 + 698],mem_3_1[0 + 699],mem_3_1[0 + 700],mem_3_1[0 + 701],mem_3_1[0 + 702],mem_3_1[0 + 703],mem_3_1[0 + 704],mem_3_1[0 + 705],mem_3_1[0 + 706],mem_3_1[0 + 707],mem_3_1[0 + 708],mem_3_1[0 + 709],mem_3_1[0 + 710],mem_3_1[0 + 711],mem_3_1[0 + 712],mem_3_1[0 + 713],mem_3_1[0 + 714],mem_3_1[0 + 715],mem_3_1[0 + 716],mem_3_1[0 + 717],mem_3_1[0 + 718],mem_3_1[0 + 719],mem_3_1[0 + 720],mem_3_1[0 + 721],mem_3_1[0 + 722],mem_3_1[0 + 723],mem_3_1[0 + 724],mem_3_1[0 + 725],mem_3_1[0 + 726],mem_3_1[0 + 727],mem_3_1[0 + 728],mem_3_1[0 + 729],mem_3_1[0 + 730],mem_3_1[0 + 731],mem_3_1[0 + 732],mem_3_1[0 + 733],mem_3_1[0 + 734],mem_3_1[0 + 735],mem_3_1[0 + 736],mem_3_1[0 + 737],mem_3_1[0 + 738],mem_3_1[0 + 739],mem_3_1[0 + 740],mem_3_1[0 + 741],mem_3_1[0 + 742],mem_3_1[0 + 743],mem_3_1[0 + 744],mem_3_1[0 + 745],mem_3_1[0 + 746],mem_3_1[0 + 747],mem_3_1[0 + 748],mem_3_1[0 + 749],mem_3_1[0 + 750],mem_3_1[0 + 751],mem_3_1[0 + 752],mem_3_1[0 + 753],mem_3_1[0 + 754],mem_3_1[0 + 755],mem_3_1[0 + 756],mem_3_1[0 + 757],mem_3_1[0 + 758],mem_3_1[0 + 759],mem_3_1[0 + 760],mem_3_1[0 + 761],mem_3_1[0 + 762],mem_3_1[0 + 763],mem_3_1[0 + 764],mem_3_1[0 + 765],mem_3_1[0 + 766],mem_3_1[0 + 767],mem_3_1[0 + 768],mem_3_1[0 + 769],mem_3_1[0 + 770],mem_3_1[0 + 771],mem_3_1[0 + 772],mem_3_1[0 + 773],mem_3_1[0 + 774],mem_3_1[0 + 775],mem_3_1[0 + 776],mem_3_1[0 + 777],mem_3_1[0 + 778],mem_3_1[0 + 779],mem_3_1[0 + 780],mem_3_1[0 + 781],mem_3_1[0 + 782],mem_3_1[0 + 783],mem_3_1[0 + 784],mem_3_1[0 + 785],mem_3_1[0 + 786],mem_3_1[0 + 787],mem_3_1[0 + 788],mem_3_1[0 + 789],mem_3_1[0 + 790],mem_3_1[0 + 791],mem_3_1[0 + 792],mem_3_1[0 + 793],mem_3_1[0 + 794],mem_3_1[0 + 795],mem_3_1[0 + 796],mem_3_1[0 + 797],mem_3_1[0 + 798],mem_3_1[0 + 799],mem_3_1[0 + 800],mem_3_1[0 + 801],mem_3_1[0 + 802],mem_3_1[0 + 803],mem_3_1[0 + 804],mem_3_1[0 + 805],mem_3_1[0 + 806],mem_3_1[0 + 807],mem_3_1[0 + 808],mem_3_1[0 + 809],mem_3_1[0 + 810],mem_3_1[0 + 811],mem_3_1[0 + 812],mem_3_1[0 + 813],mem_3_1[0 + 814],mem_3_1[0 + 815],mem_3_1[0 + 816],mem_3_1[0 + 817],mem_3_1[0 + 818],mem_3_1[0 + 819],mem_3_1[0 + 820],mem_3_1[0 + 821],mem_3_1[0 + 822],mem_3_1[0 + 823],mem_3_1[0 + 824],mem_3_1[0 + 825],mem_3_1[0 + 826],mem_3_1[0 + 827],mem_3_1[0 + 828],mem_3_1[0 + 829],mem_3_1[0 + 830],mem_3_1[0 + 831],mem_3_1[0 + 832],mem_3_1[0 + 833],mem_3_1[0 + 834],mem_3_1[0 + 835],mem_3_1[0 + 836],mem_3_1[0 + 837],mem_3_1[0 + 838],mem_3_1[0 + 839],mem_3_1[0 + 840],mem_3_1[0 + 841],mem_3_1[0 + 842],mem_3_1[0 + 843],mem_3_1[0 + 844],mem_3_1[0 + 845],mem_3_1[0 + 846],mem_3_1[0 + 847],mem_3_1[0 + 848],mem_3_1[0 + 849],mem_3_1[0 + 850],mem_3_1[0 + 851],mem_3_1[0 + 852],mem_3_1[0 + 853],mem_3_1[0 + 854],mem_3_1[0 + 855],mem_3_1[0 + 856],mem_3_1[0 + 857],mem_3_1[0 + 858],mem_3_1[0 + 859],mem_3_1[0 + 860],mem_3_1[0 + 861],mem_3_1[0 + 862],mem_3_1[0 + 863],mem_3_1[0 + 864],mem_3_1[0 + 865],mem_3_1[0 + 866],mem_3_1[0 + 867],mem_3_1[0 + 868],mem_3_1[0 + 869],mem_3_1[0 + 870],mem_3_1[0 + 871],mem_3_1[0 + 872],mem_3_1[0 + 873],mem_3_1[0 + 874],mem_3_1[0 + 875],mem_3_1[0 + 876],mem_3_1[0 + 877],mem_3_1[0 + 878],mem_3_1[0 + 879],mem_3_1[0 + 880],mem_3_1[0 + 881],mem_3_1[0 + 882],mem_3_1[0 + 883],mem_3_1[0 + 884],mem_3_1[0 + 885],mem_3_1[0 + 886],mem_3_1[0 + 887],mem_3_1[0 + 888],mem_3_1[0 + 889],mem_3_1[0 + 890],mem_3_1[0 + 891],mem_3_1[0 + 892],mem_3_1[0 + 893],mem_3_1[0 + 894],mem_3_1[0 + 895],mem_3_1[0 + 896],mem_3_1[0 + 897],mem_3_1[0 + 898],mem_3_1[0 + 899],mem_3_1[0 + 900],mem_3_1[0 + 901],mem_3_1[0 + 902],mem_3_1[0 + 903],mem_3_1[0 + 904],mem_3_1[0 + 905],mem_3_1[0 + 906],mem_3_1[0 + 907],mem_3_1[0 + 908],mem_3_1[0 + 909],mem_3_1[0 + 910],mem_3_1[0 + 911],mem_3_1[0 + 912],mem_3_1[0 + 913],mem_3_1[0 + 914],mem_3_1[0 + 915],mem_3_1[0 + 916],mem_3_1[0 + 917],mem_3_1[0 + 918],mem_3_1[0 + 919],mem_3_1[0 + 920],mem_3_1[0 + 921],mem_3_1[0 + 922],mem_3_1[0 + 923],mem_3_1[0 + 924],mem_3_1[0 + 925],mem_3_1[0 + 926],mem_3_1[0 + 927],mem_3_1[0 + 928],mem_3_1[0 + 929],mem_3_1[0 + 930],mem_3_1[0 + 931],mem_3_1[0 + 932],mem_3_1[0 + 933],mem_3_1[0 + 934],mem_3_1[0 + 935],mem_3_1[0 + 936],mem_3_1[0 + 937],mem_3_1[0 + 938],mem_3_1[0 + 939],mem_3_1[0 + 940],mem_3_1[0 + 941],mem_3_1[0 + 942],mem_3_1[0 + 943],mem_3_1[0 + 944],mem_3_1[0 + 945],mem_3_1[0 + 946],mem_3_1[0 + 947],mem_3_1[0 + 948],mem_3_1[0 + 949],mem_3_1[0 + 950],mem_3_1[0 + 951],mem_3_1[0 + 952],mem_3_1[0 + 953],mem_3_1[0 + 954],mem_3_1[0 + 955],mem_3_1[0 + 956],mem_3_1[0 + 957],mem_3_1[0 + 958],mem_3_1[0 + 959],mem_3_1[0 + 960],mem_3_1[0 + 961],mem_3_1[0 + 962],mem_3_1[0 + 963],mem_3_1[0 + 964],mem_3_1[0 + 965],mem_3_1[0 + 966],mem_3_1[0 + 967],mem_3_1[0 + 968],mem_3_1[0 + 969],mem_3_1[0 + 970],mem_3_1[0 + 971],mem_3_1[0 + 972],mem_3_1[0 + 973],mem_3_1[0 + 974],mem_3_1[0 + 975],mem_3_1[0 + 976],mem_3_1[0 + 977],mem_3_1[0 + 978],mem_3_1[0 + 979],mem_3_1[0 + 980],mem_3_1[0 + 981],mem_3_1[0 + 982],mem_3_1[0 + 983],mem_3_1[0 + 984],mem_3_1[0 + 985],mem_3_1[0 + 986],mem_3_1[0 + 987],mem_3_1[0 + 988],mem_3_1[0 + 989],mem_3_1[0 + 990],mem_3_1[0 + 991],mem_3_1[0 + 992],mem_3_1[0 + 993],mem_3_1[0 + 994],mem_3_1[0 + 995],mem_3_1[0 + 996],mem_3_1[0 + 997],mem_3_1[0 + 998],mem_3_1[0 + 999],mem_3_1[0 + 1000],mem_3_1[0 + 1001],mem_3_1[0 + 1002],mem_3_1[0 + 1003],mem_3_1[0 + 1004],mem_3_1[0 + 1005],mem_3_1[0 + 1006],mem_3_1[0 + 1007],mem_3_1[0 + 1008],mem_3_1[0 + 1009],mem_3_1[0 + 1010],mem_3_1[0 + 1011],mem_3_1[0 + 1012],mem_3_1[0 + 1013],mem_3_1[0 + 1014],mem_3_1[0 + 1015],mem_3_1[0 + 1016],mem_3_1[0 + 1017],mem_3_1[0 + 1018],mem_3_1[0 + 1019],mem_3_1[0 + 1020],mem_3_1[0 + 1021],mem_3_1[0 + 1022],mem_3_1[0 + 1024 - 1] };
wire [8*(1024)-1:0] mem_0_0_flat_src;
assign mem_0_0_flat_src = {mem_0_0[0 + 0],mem_0_0[0 + 1],mem_0_0[0 + 2],mem_0_0[0 + 3],mem_0_0[0 + 4],mem_0_0[0 + 5],mem_0_0[0 + 6],mem_0_0[0 + 7],mem_0_0[0 + 8],mem_0_0[0 + 9],mem_0_0[0 + 10],mem_0_0[0 + 11],mem_0_0[0 + 12],mem_0_0[0 + 13],mem_0_0[0 + 14],mem_0_0[0 + 15],mem_0_0[0 + 16],mem_0_0[0 + 17],mem_0_0[0 + 18],mem_0_0[0 + 19],mem_0_0[0 + 20],mem_0_0[0 + 21],mem_0_0[0 + 22],mem_0_0[0 + 23],mem_0_0[0 + 24],mem_0_0[0 + 25],mem_0_0[0 + 26],mem_0_0[0 + 27],mem_0_0[0 + 28],mem_0_0[0 + 29],mem_0_0[0 + 30],mem_0_0[0 + 31],mem_0_0[0 + 32],mem_0_0[0 + 33],mem_0_0[0 + 34],mem_0_0[0 + 35],mem_0_0[0 + 36],mem_0_0[0 + 37],mem_0_0[0 + 38],mem_0_0[0 + 39],mem_0_0[0 + 40],mem_0_0[0 + 41],mem_0_0[0 + 42],mem_0_0[0 + 43],mem_0_0[0 + 44],mem_0_0[0 + 45],mem_0_0[0 + 46],mem_0_0[0 + 47],mem_0_0[0 + 48],mem_0_0[0 + 49],mem_0_0[0 + 50],mem_0_0[0 + 51],mem_0_0[0 + 52],mem_0_0[0 + 53],mem_0_0[0 + 54],mem_0_0[0 + 55],mem_0_0[0 + 56],mem_0_0[0 + 57],mem_0_0[0 + 58],mem_0_0[0 + 59],mem_0_0[0 + 60],mem_0_0[0 + 61],mem_0_0[0 + 62],mem_0_0[0 + 63],mem_0_0[0 + 64],mem_0_0[0 + 65],mem_0_0[0 + 66],mem_0_0[0 + 67],mem_0_0[0 + 68],mem_0_0[0 + 69],mem_0_0[0 + 70],mem_0_0[0 + 71],mem_0_0[0 + 72],mem_0_0[0 + 73],mem_0_0[0 + 74],mem_0_0[0 + 75],mem_0_0[0 + 76],mem_0_0[0 + 77],mem_0_0[0 + 78],mem_0_0[0 + 79],mem_0_0[0 + 80],mem_0_0[0 + 81],mem_0_0[0 + 82],mem_0_0[0 + 83],mem_0_0[0 + 84],mem_0_0[0 + 85],mem_0_0[0 + 86],mem_0_0[0 + 87],mem_0_0[0 + 88],mem_0_0[0 + 89],mem_0_0[0 + 90],mem_0_0[0 + 91],mem_0_0[0 + 92],mem_0_0[0 + 93],mem_0_0[0 + 94],mem_0_0[0 + 95],mem_0_0[0 + 96],mem_0_0[0 + 97],mem_0_0[0 + 98],mem_0_0[0 + 99],mem_0_0[0 + 100],mem_0_0[0 + 101],mem_0_0[0 + 102],mem_0_0[0 + 103],mem_0_0[0 + 104],mem_0_0[0 + 105],mem_0_0[0 + 106],mem_0_0[0 + 107],mem_0_0[0 + 108],mem_0_0[0 + 109],mem_0_0[0 + 110],mem_0_0[0 + 111],mem_0_0[0 + 112],mem_0_0[0 + 113],mem_0_0[0 + 114],mem_0_0[0 + 115],mem_0_0[0 + 116],mem_0_0[0 + 117],mem_0_0[0 + 118],mem_0_0[0 + 119],mem_0_0[0 + 120],mem_0_0[0 + 121],mem_0_0[0 + 122],mem_0_0[0 + 123],mem_0_0[0 + 124],mem_0_0[0 + 125],mem_0_0[0 + 126],mem_0_0[0 + 127],mem_0_0[0 + 128],mem_0_0[0 + 129],mem_0_0[0 + 130],mem_0_0[0 + 131],mem_0_0[0 + 132],mem_0_0[0 + 133],mem_0_0[0 + 134],mem_0_0[0 + 135],mem_0_0[0 + 136],mem_0_0[0 + 137],mem_0_0[0 + 138],mem_0_0[0 + 139],mem_0_0[0 + 140],mem_0_0[0 + 141],mem_0_0[0 + 142],mem_0_0[0 + 143],mem_0_0[0 + 144],mem_0_0[0 + 145],mem_0_0[0 + 146],mem_0_0[0 + 147],mem_0_0[0 + 148],mem_0_0[0 + 149],mem_0_0[0 + 150],mem_0_0[0 + 151],mem_0_0[0 + 152],mem_0_0[0 + 153],mem_0_0[0 + 154],mem_0_0[0 + 155],mem_0_0[0 + 156],mem_0_0[0 + 157],mem_0_0[0 + 158],mem_0_0[0 + 159],mem_0_0[0 + 160],mem_0_0[0 + 161],mem_0_0[0 + 162],mem_0_0[0 + 163],mem_0_0[0 + 164],mem_0_0[0 + 165],mem_0_0[0 + 166],mem_0_0[0 + 167],mem_0_0[0 + 168],mem_0_0[0 + 169],mem_0_0[0 + 170],mem_0_0[0 + 171],mem_0_0[0 + 172],mem_0_0[0 + 173],mem_0_0[0 + 174],mem_0_0[0 + 175],mem_0_0[0 + 176],mem_0_0[0 + 177],mem_0_0[0 + 178],mem_0_0[0 + 179],mem_0_0[0 + 180],mem_0_0[0 + 181],mem_0_0[0 + 182],mem_0_0[0 + 183],mem_0_0[0 + 184],mem_0_0[0 + 185],mem_0_0[0 + 186],mem_0_0[0 + 187],mem_0_0[0 + 188],mem_0_0[0 + 189],mem_0_0[0 + 190],mem_0_0[0 + 191],mem_0_0[0 + 192],mem_0_0[0 + 193],mem_0_0[0 + 194],mem_0_0[0 + 195],mem_0_0[0 + 196],mem_0_0[0 + 197],mem_0_0[0 + 198],mem_0_0[0 + 199],mem_0_0[0 + 200],mem_0_0[0 + 201],mem_0_0[0 + 202],mem_0_0[0 + 203],mem_0_0[0 + 204],mem_0_0[0 + 205],mem_0_0[0 + 206],mem_0_0[0 + 207],mem_0_0[0 + 208],mem_0_0[0 + 209],mem_0_0[0 + 210],mem_0_0[0 + 211],mem_0_0[0 + 212],mem_0_0[0 + 213],mem_0_0[0 + 214],mem_0_0[0 + 215],mem_0_0[0 + 216],mem_0_0[0 + 217],mem_0_0[0 + 218],mem_0_0[0 + 219],mem_0_0[0 + 220],mem_0_0[0 + 221],mem_0_0[0 + 222],mem_0_0[0 + 223],mem_0_0[0 + 224],mem_0_0[0 + 225],mem_0_0[0 + 226],mem_0_0[0 + 227],mem_0_0[0 + 228],mem_0_0[0 + 229],mem_0_0[0 + 230],mem_0_0[0 + 231],mem_0_0[0 + 232],mem_0_0[0 + 233],mem_0_0[0 + 234],mem_0_0[0 + 235],mem_0_0[0 + 236],mem_0_0[0 + 237],mem_0_0[0 + 238],mem_0_0[0 + 239],mem_0_0[0 + 240],mem_0_0[0 + 241],mem_0_0[0 + 242],mem_0_0[0 + 243],mem_0_0[0 + 244],mem_0_0[0 + 245],mem_0_0[0 + 246],mem_0_0[0 + 247],mem_0_0[0 + 248],mem_0_0[0 + 249],mem_0_0[0 + 250],mem_0_0[0 + 251],mem_0_0[0 + 252],mem_0_0[0 + 253],mem_0_0[0 + 254],mem_0_0[0 + 255],mem_0_0[0 + 256],mem_0_0[0 + 257],mem_0_0[0 + 258],mem_0_0[0 + 259],mem_0_0[0 + 260],mem_0_0[0 + 261],mem_0_0[0 + 262],mem_0_0[0 + 263],mem_0_0[0 + 264],mem_0_0[0 + 265],mem_0_0[0 + 266],mem_0_0[0 + 267],mem_0_0[0 + 268],mem_0_0[0 + 269],mem_0_0[0 + 270],mem_0_0[0 + 271],mem_0_0[0 + 272],mem_0_0[0 + 273],mem_0_0[0 + 274],mem_0_0[0 + 275],mem_0_0[0 + 276],mem_0_0[0 + 277],mem_0_0[0 + 278],mem_0_0[0 + 279],mem_0_0[0 + 280],mem_0_0[0 + 281],mem_0_0[0 + 282],mem_0_0[0 + 283],mem_0_0[0 + 284],mem_0_0[0 + 285],mem_0_0[0 + 286],mem_0_0[0 + 287],mem_0_0[0 + 288],mem_0_0[0 + 289],mem_0_0[0 + 290],mem_0_0[0 + 291],mem_0_0[0 + 292],mem_0_0[0 + 293],mem_0_0[0 + 294],mem_0_0[0 + 295],mem_0_0[0 + 296],mem_0_0[0 + 297],mem_0_0[0 + 298],mem_0_0[0 + 299],mem_0_0[0 + 300],mem_0_0[0 + 301],mem_0_0[0 + 302],mem_0_0[0 + 303],mem_0_0[0 + 304],mem_0_0[0 + 305],mem_0_0[0 + 306],mem_0_0[0 + 307],mem_0_0[0 + 308],mem_0_0[0 + 309],mem_0_0[0 + 310],mem_0_0[0 + 311],mem_0_0[0 + 312],mem_0_0[0 + 313],mem_0_0[0 + 314],mem_0_0[0 + 315],mem_0_0[0 + 316],mem_0_0[0 + 317],mem_0_0[0 + 318],mem_0_0[0 + 319],mem_0_0[0 + 320],mem_0_0[0 + 321],mem_0_0[0 + 322],mem_0_0[0 + 323],mem_0_0[0 + 324],mem_0_0[0 + 325],mem_0_0[0 + 326],mem_0_0[0 + 327],mem_0_0[0 + 328],mem_0_0[0 + 329],mem_0_0[0 + 330],mem_0_0[0 + 331],mem_0_0[0 + 332],mem_0_0[0 + 333],mem_0_0[0 + 334],mem_0_0[0 + 335],mem_0_0[0 + 336],mem_0_0[0 + 337],mem_0_0[0 + 338],mem_0_0[0 + 339],mem_0_0[0 + 340],mem_0_0[0 + 341],mem_0_0[0 + 342],mem_0_0[0 + 343],mem_0_0[0 + 344],mem_0_0[0 + 345],mem_0_0[0 + 346],mem_0_0[0 + 347],mem_0_0[0 + 348],mem_0_0[0 + 349],mem_0_0[0 + 350],mem_0_0[0 + 351],mem_0_0[0 + 352],mem_0_0[0 + 353],mem_0_0[0 + 354],mem_0_0[0 + 355],mem_0_0[0 + 356],mem_0_0[0 + 357],mem_0_0[0 + 358],mem_0_0[0 + 359],mem_0_0[0 + 360],mem_0_0[0 + 361],mem_0_0[0 + 362],mem_0_0[0 + 363],mem_0_0[0 + 364],mem_0_0[0 + 365],mem_0_0[0 + 366],mem_0_0[0 + 367],mem_0_0[0 + 368],mem_0_0[0 + 369],mem_0_0[0 + 370],mem_0_0[0 + 371],mem_0_0[0 + 372],mem_0_0[0 + 373],mem_0_0[0 + 374],mem_0_0[0 + 375],mem_0_0[0 + 376],mem_0_0[0 + 377],mem_0_0[0 + 378],mem_0_0[0 + 379],mem_0_0[0 + 380],mem_0_0[0 + 381],mem_0_0[0 + 382],mem_0_0[0 + 383],mem_0_0[0 + 384],mem_0_0[0 + 385],mem_0_0[0 + 386],mem_0_0[0 + 387],mem_0_0[0 + 388],mem_0_0[0 + 389],mem_0_0[0 + 390],mem_0_0[0 + 391],mem_0_0[0 + 392],mem_0_0[0 + 393],mem_0_0[0 + 394],mem_0_0[0 + 395],mem_0_0[0 + 396],mem_0_0[0 + 397],mem_0_0[0 + 398],mem_0_0[0 + 399],mem_0_0[0 + 400],mem_0_0[0 + 401],mem_0_0[0 + 402],mem_0_0[0 + 403],mem_0_0[0 + 404],mem_0_0[0 + 405],mem_0_0[0 + 406],mem_0_0[0 + 407],mem_0_0[0 + 408],mem_0_0[0 + 409],mem_0_0[0 + 410],mem_0_0[0 + 411],mem_0_0[0 + 412],mem_0_0[0 + 413],mem_0_0[0 + 414],mem_0_0[0 + 415],mem_0_0[0 + 416],mem_0_0[0 + 417],mem_0_0[0 + 418],mem_0_0[0 + 419],mem_0_0[0 + 420],mem_0_0[0 + 421],mem_0_0[0 + 422],mem_0_0[0 + 423],mem_0_0[0 + 424],mem_0_0[0 + 425],mem_0_0[0 + 426],mem_0_0[0 + 427],mem_0_0[0 + 428],mem_0_0[0 + 429],mem_0_0[0 + 430],mem_0_0[0 + 431],mem_0_0[0 + 432],mem_0_0[0 + 433],mem_0_0[0 + 434],mem_0_0[0 + 435],mem_0_0[0 + 436],mem_0_0[0 + 437],mem_0_0[0 + 438],mem_0_0[0 + 439],mem_0_0[0 + 440],mem_0_0[0 + 441],mem_0_0[0 + 442],mem_0_0[0 + 443],mem_0_0[0 + 444],mem_0_0[0 + 445],mem_0_0[0 + 446],mem_0_0[0 + 447],mem_0_0[0 + 448],mem_0_0[0 + 449],mem_0_0[0 + 450],mem_0_0[0 + 451],mem_0_0[0 + 452],mem_0_0[0 + 453],mem_0_0[0 + 454],mem_0_0[0 + 455],mem_0_0[0 + 456],mem_0_0[0 + 457],mem_0_0[0 + 458],mem_0_0[0 + 459],mem_0_0[0 + 460],mem_0_0[0 + 461],mem_0_0[0 + 462],mem_0_0[0 + 463],mem_0_0[0 + 464],mem_0_0[0 + 465],mem_0_0[0 + 466],mem_0_0[0 + 467],mem_0_0[0 + 468],mem_0_0[0 + 469],mem_0_0[0 + 470],mem_0_0[0 + 471],mem_0_0[0 + 472],mem_0_0[0 + 473],mem_0_0[0 + 474],mem_0_0[0 + 475],mem_0_0[0 + 476],mem_0_0[0 + 477],mem_0_0[0 + 478],mem_0_0[0 + 479],mem_0_0[0 + 480],mem_0_0[0 + 481],mem_0_0[0 + 482],mem_0_0[0 + 483],mem_0_0[0 + 484],mem_0_0[0 + 485],mem_0_0[0 + 486],mem_0_0[0 + 487],mem_0_0[0 + 488],mem_0_0[0 + 489],mem_0_0[0 + 490],mem_0_0[0 + 491],mem_0_0[0 + 492],mem_0_0[0 + 493],mem_0_0[0 + 494],mem_0_0[0 + 495],mem_0_0[0 + 496],mem_0_0[0 + 497],mem_0_0[0 + 498],mem_0_0[0 + 499],mem_0_0[0 + 500],mem_0_0[0 + 501],mem_0_0[0 + 502],mem_0_0[0 + 503],mem_0_0[0 + 504],mem_0_0[0 + 505],mem_0_0[0 + 506],mem_0_0[0 + 507],mem_0_0[0 + 508],mem_0_0[0 + 509],mem_0_0[0 + 510],mem_0_0[0 + 511],mem_0_0[0 + 512],mem_0_0[0 + 513],mem_0_0[0 + 514],mem_0_0[0 + 515],mem_0_0[0 + 516],mem_0_0[0 + 517],mem_0_0[0 + 518],mem_0_0[0 + 519],mem_0_0[0 + 520],mem_0_0[0 + 521],mem_0_0[0 + 522],mem_0_0[0 + 523],mem_0_0[0 + 524],mem_0_0[0 + 525],mem_0_0[0 + 526],mem_0_0[0 + 527],mem_0_0[0 + 528],mem_0_0[0 + 529],mem_0_0[0 + 530],mem_0_0[0 + 531],mem_0_0[0 + 532],mem_0_0[0 + 533],mem_0_0[0 + 534],mem_0_0[0 + 535],mem_0_0[0 + 536],mem_0_0[0 + 537],mem_0_0[0 + 538],mem_0_0[0 + 539],mem_0_0[0 + 540],mem_0_0[0 + 541],mem_0_0[0 + 542],mem_0_0[0 + 543],mem_0_0[0 + 544],mem_0_0[0 + 545],mem_0_0[0 + 546],mem_0_0[0 + 547],mem_0_0[0 + 548],mem_0_0[0 + 549],mem_0_0[0 + 550],mem_0_0[0 + 551],mem_0_0[0 + 552],mem_0_0[0 + 553],mem_0_0[0 + 554],mem_0_0[0 + 555],mem_0_0[0 + 556],mem_0_0[0 + 557],mem_0_0[0 + 558],mem_0_0[0 + 559],mem_0_0[0 + 560],mem_0_0[0 + 561],mem_0_0[0 + 562],mem_0_0[0 + 563],mem_0_0[0 + 564],mem_0_0[0 + 565],mem_0_0[0 + 566],mem_0_0[0 + 567],mem_0_0[0 + 568],mem_0_0[0 + 569],mem_0_0[0 + 570],mem_0_0[0 + 571],mem_0_0[0 + 572],mem_0_0[0 + 573],mem_0_0[0 + 574],mem_0_0[0 + 575],mem_0_0[0 + 576],mem_0_0[0 + 577],mem_0_0[0 + 578],mem_0_0[0 + 579],mem_0_0[0 + 580],mem_0_0[0 + 581],mem_0_0[0 + 582],mem_0_0[0 + 583],mem_0_0[0 + 584],mem_0_0[0 + 585],mem_0_0[0 + 586],mem_0_0[0 + 587],mem_0_0[0 + 588],mem_0_0[0 + 589],mem_0_0[0 + 590],mem_0_0[0 + 591],mem_0_0[0 + 592],mem_0_0[0 + 593],mem_0_0[0 + 594],mem_0_0[0 + 595],mem_0_0[0 + 596],mem_0_0[0 + 597],mem_0_0[0 + 598],mem_0_0[0 + 599],mem_0_0[0 + 600],mem_0_0[0 + 601],mem_0_0[0 + 602],mem_0_0[0 + 603],mem_0_0[0 + 604],mem_0_0[0 + 605],mem_0_0[0 + 606],mem_0_0[0 + 607],mem_0_0[0 + 608],mem_0_0[0 + 609],mem_0_0[0 + 610],mem_0_0[0 + 611],mem_0_0[0 + 612],mem_0_0[0 + 613],mem_0_0[0 + 614],mem_0_0[0 + 615],mem_0_0[0 + 616],mem_0_0[0 + 617],mem_0_0[0 + 618],mem_0_0[0 + 619],mem_0_0[0 + 620],mem_0_0[0 + 621],mem_0_0[0 + 622],mem_0_0[0 + 623],mem_0_0[0 + 624],mem_0_0[0 + 625],mem_0_0[0 + 626],mem_0_0[0 + 627],mem_0_0[0 + 628],mem_0_0[0 + 629],mem_0_0[0 + 630],mem_0_0[0 + 631],mem_0_0[0 + 632],mem_0_0[0 + 633],mem_0_0[0 + 634],mem_0_0[0 + 635],mem_0_0[0 + 636],mem_0_0[0 + 637],mem_0_0[0 + 638],mem_0_0[0 + 639],mem_0_0[0 + 640],mem_0_0[0 + 641],mem_0_0[0 + 642],mem_0_0[0 + 643],mem_0_0[0 + 644],mem_0_0[0 + 645],mem_0_0[0 + 646],mem_0_0[0 + 647],mem_0_0[0 + 648],mem_0_0[0 + 649],mem_0_0[0 + 650],mem_0_0[0 + 651],mem_0_0[0 + 652],mem_0_0[0 + 653],mem_0_0[0 + 654],mem_0_0[0 + 655],mem_0_0[0 + 656],mem_0_0[0 + 657],mem_0_0[0 + 658],mem_0_0[0 + 659],mem_0_0[0 + 660],mem_0_0[0 + 661],mem_0_0[0 + 662],mem_0_0[0 + 663],mem_0_0[0 + 664],mem_0_0[0 + 665],mem_0_0[0 + 666],mem_0_0[0 + 667],mem_0_0[0 + 668],mem_0_0[0 + 669],mem_0_0[0 + 670],mem_0_0[0 + 671],mem_0_0[0 + 672],mem_0_0[0 + 673],mem_0_0[0 + 674],mem_0_0[0 + 675],mem_0_0[0 + 676],mem_0_0[0 + 677],mem_0_0[0 + 678],mem_0_0[0 + 679],mem_0_0[0 + 680],mem_0_0[0 + 681],mem_0_0[0 + 682],mem_0_0[0 + 683],mem_0_0[0 + 684],mem_0_0[0 + 685],mem_0_0[0 + 686],mem_0_0[0 + 687],mem_0_0[0 + 688],mem_0_0[0 + 689],mem_0_0[0 + 690],mem_0_0[0 + 691],mem_0_0[0 + 692],mem_0_0[0 + 693],mem_0_0[0 + 694],mem_0_0[0 + 695],mem_0_0[0 + 696],mem_0_0[0 + 697],mem_0_0[0 + 698],mem_0_0[0 + 699],mem_0_0[0 + 700],mem_0_0[0 + 701],mem_0_0[0 + 702],mem_0_0[0 + 703],mem_0_0[0 + 704],mem_0_0[0 + 705],mem_0_0[0 + 706],mem_0_0[0 + 707],mem_0_0[0 + 708],mem_0_0[0 + 709],mem_0_0[0 + 710],mem_0_0[0 + 711],mem_0_0[0 + 712],mem_0_0[0 + 713],mem_0_0[0 + 714],mem_0_0[0 + 715],mem_0_0[0 + 716],mem_0_0[0 + 717],mem_0_0[0 + 718],mem_0_0[0 + 719],mem_0_0[0 + 720],mem_0_0[0 + 721],mem_0_0[0 + 722],mem_0_0[0 + 723],mem_0_0[0 + 724],mem_0_0[0 + 725],mem_0_0[0 + 726],mem_0_0[0 + 727],mem_0_0[0 + 728],mem_0_0[0 + 729],mem_0_0[0 + 730],mem_0_0[0 + 731],mem_0_0[0 + 732],mem_0_0[0 + 733],mem_0_0[0 + 734],mem_0_0[0 + 735],mem_0_0[0 + 736],mem_0_0[0 + 737],mem_0_0[0 + 738],mem_0_0[0 + 739],mem_0_0[0 + 740],mem_0_0[0 + 741],mem_0_0[0 + 742],mem_0_0[0 + 743],mem_0_0[0 + 744],mem_0_0[0 + 745],mem_0_0[0 + 746],mem_0_0[0 + 747],mem_0_0[0 + 748],mem_0_0[0 + 749],mem_0_0[0 + 750],mem_0_0[0 + 751],mem_0_0[0 + 752],mem_0_0[0 + 753],mem_0_0[0 + 754],mem_0_0[0 + 755],mem_0_0[0 + 756],mem_0_0[0 + 757],mem_0_0[0 + 758],mem_0_0[0 + 759],mem_0_0[0 + 760],mem_0_0[0 + 761],mem_0_0[0 + 762],mem_0_0[0 + 763],mem_0_0[0 + 764],mem_0_0[0 + 765],mem_0_0[0 + 766],mem_0_0[0 + 767],mem_0_0[0 + 768],mem_0_0[0 + 769],mem_0_0[0 + 770],mem_0_0[0 + 771],mem_0_0[0 + 772],mem_0_0[0 + 773],mem_0_0[0 + 774],mem_0_0[0 + 775],mem_0_0[0 + 776],mem_0_0[0 + 777],mem_0_0[0 + 778],mem_0_0[0 + 779],mem_0_0[0 + 780],mem_0_0[0 + 781],mem_0_0[0 + 782],mem_0_0[0 + 783],mem_0_0[0 + 784],mem_0_0[0 + 785],mem_0_0[0 + 786],mem_0_0[0 + 787],mem_0_0[0 + 788],mem_0_0[0 + 789],mem_0_0[0 + 790],mem_0_0[0 + 791],mem_0_0[0 + 792],mem_0_0[0 + 793],mem_0_0[0 + 794],mem_0_0[0 + 795],mem_0_0[0 + 796],mem_0_0[0 + 797],mem_0_0[0 + 798],mem_0_0[0 + 799],mem_0_0[0 + 800],mem_0_0[0 + 801],mem_0_0[0 + 802],mem_0_0[0 + 803],mem_0_0[0 + 804],mem_0_0[0 + 805],mem_0_0[0 + 806],mem_0_0[0 + 807],mem_0_0[0 + 808],mem_0_0[0 + 809],mem_0_0[0 + 810],mem_0_0[0 + 811],mem_0_0[0 + 812],mem_0_0[0 + 813],mem_0_0[0 + 814],mem_0_0[0 + 815],mem_0_0[0 + 816],mem_0_0[0 + 817],mem_0_0[0 + 818],mem_0_0[0 + 819],mem_0_0[0 + 820],mem_0_0[0 + 821],mem_0_0[0 + 822],mem_0_0[0 + 823],mem_0_0[0 + 824],mem_0_0[0 + 825],mem_0_0[0 + 826],mem_0_0[0 + 827],mem_0_0[0 + 828],mem_0_0[0 + 829],mem_0_0[0 + 830],mem_0_0[0 + 831],mem_0_0[0 + 832],mem_0_0[0 + 833],mem_0_0[0 + 834],mem_0_0[0 + 835],mem_0_0[0 + 836],mem_0_0[0 + 837],mem_0_0[0 + 838],mem_0_0[0 + 839],mem_0_0[0 + 840],mem_0_0[0 + 841],mem_0_0[0 + 842],mem_0_0[0 + 843],mem_0_0[0 + 844],mem_0_0[0 + 845],mem_0_0[0 + 846],mem_0_0[0 + 847],mem_0_0[0 + 848],mem_0_0[0 + 849],mem_0_0[0 + 850],mem_0_0[0 + 851],mem_0_0[0 + 852],mem_0_0[0 + 853],mem_0_0[0 + 854],mem_0_0[0 + 855],mem_0_0[0 + 856],mem_0_0[0 + 857],mem_0_0[0 + 858],mem_0_0[0 + 859],mem_0_0[0 + 860],mem_0_0[0 + 861],mem_0_0[0 + 862],mem_0_0[0 + 863],mem_0_0[0 + 864],mem_0_0[0 + 865],mem_0_0[0 + 866],mem_0_0[0 + 867],mem_0_0[0 + 868],mem_0_0[0 + 869],mem_0_0[0 + 870],mem_0_0[0 + 871],mem_0_0[0 + 872],mem_0_0[0 + 873],mem_0_0[0 + 874],mem_0_0[0 + 875],mem_0_0[0 + 876],mem_0_0[0 + 877],mem_0_0[0 + 878],mem_0_0[0 + 879],mem_0_0[0 + 880],mem_0_0[0 + 881],mem_0_0[0 + 882],mem_0_0[0 + 883],mem_0_0[0 + 884],mem_0_0[0 + 885],mem_0_0[0 + 886],mem_0_0[0 + 887],mem_0_0[0 + 888],mem_0_0[0 + 889],mem_0_0[0 + 890],mem_0_0[0 + 891],mem_0_0[0 + 892],mem_0_0[0 + 893],mem_0_0[0 + 894],mem_0_0[0 + 895],mem_0_0[0 + 896],mem_0_0[0 + 897],mem_0_0[0 + 898],mem_0_0[0 + 899],mem_0_0[0 + 900],mem_0_0[0 + 901],mem_0_0[0 + 902],mem_0_0[0 + 903],mem_0_0[0 + 904],mem_0_0[0 + 905],mem_0_0[0 + 906],mem_0_0[0 + 907],mem_0_0[0 + 908],mem_0_0[0 + 909],mem_0_0[0 + 910],mem_0_0[0 + 911],mem_0_0[0 + 912],mem_0_0[0 + 913],mem_0_0[0 + 914],mem_0_0[0 + 915],mem_0_0[0 + 916],mem_0_0[0 + 917],mem_0_0[0 + 918],mem_0_0[0 + 919],mem_0_0[0 + 920],mem_0_0[0 + 921],mem_0_0[0 + 922],mem_0_0[0 + 923],mem_0_0[0 + 924],mem_0_0[0 + 925],mem_0_0[0 + 926],mem_0_0[0 + 927],mem_0_0[0 + 928],mem_0_0[0 + 929],mem_0_0[0 + 930],mem_0_0[0 + 931],mem_0_0[0 + 932],mem_0_0[0 + 933],mem_0_0[0 + 934],mem_0_0[0 + 935],mem_0_0[0 + 936],mem_0_0[0 + 937],mem_0_0[0 + 938],mem_0_0[0 + 939],mem_0_0[0 + 940],mem_0_0[0 + 941],mem_0_0[0 + 942],mem_0_0[0 + 943],mem_0_0[0 + 944],mem_0_0[0 + 945],mem_0_0[0 + 946],mem_0_0[0 + 947],mem_0_0[0 + 948],mem_0_0[0 + 949],mem_0_0[0 + 950],mem_0_0[0 + 951],mem_0_0[0 + 952],mem_0_0[0 + 953],mem_0_0[0 + 954],mem_0_0[0 + 955],mem_0_0[0 + 956],mem_0_0[0 + 957],mem_0_0[0 + 958],mem_0_0[0 + 959],mem_0_0[0 + 960],mem_0_0[0 + 961],mem_0_0[0 + 962],mem_0_0[0 + 963],mem_0_0[0 + 964],mem_0_0[0 + 965],mem_0_0[0 + 966],mem_0_0[0 + 967],mem_0_0[0 + 968],mem_0_0[0 + 969],mem_0_0[0 + 970],mem_0_0[0 + 971],mem_0_0[0 + 972],mem_0_0[0 + 973],mem_0_0[0 + 974],mem_0_0[0 + 975],mem_0_0[0 + 976],mem_0_0[0 + 977],mem_0_0[0 + 978],mem_0_0[0 + 979],mem_0_0[0 + 980],mem_0_0[0 + 981],mem_0_0[0 + 982],mem_0_0[0 + 983],mem_0_0[0 + 984],mem_0_0[0 + 985],mem_0_0[0 + 986],mem_0_0[0 + 987],mem_0_0[0 + 988],mem_0_0[0 + 989],mem_0_0[0 + 990],mem_0_0[0 + 991],mem_0_0[0 + 992],mem_0_0[0 + 993],mem_0_0[0 + 994],mem_0_0[0 + 995],mem_0_0[0 + 996],mem_0_0[0 + 997],mem_0_0[0 + 998],mem_0_0[0 + 999],mem_0_0[0 + 1000],mem_0_0[0 + 1001],mem_0_0[0 + 1002],mem_0_0[0 + 1003],mem_0_0[0 + 1004],mem_0_0[0 + 1005],mem_0_0[0 + 1006],mem_0_0[0 + 1007],mem_0_0[0 + 1008],mem_0_0[0 + 1009],mem_0_0[0 + 1010],mem_0_0[0 + 1011],mem_0_0[0 + 1012],mem_0_0[0 + 1013],mem_0_0[0 + 1014],mem_0_0[0 + 1015],mem_0_0[0 + 1016],mem_0_0[0 + 1017],mem_0_0[0 + 1018],mem_0_0[0 + 1019],mem_0_0[0 + 1020],mem_0_0[0 + 1021],mem_0_0[0 + 1022],mem_0_0[0 + 1024 - 1] };
wire [8*(1024)-1:0] mem_1_0_flat_src;
assign mem_1_0_flat_src = {mem_1_0[0 + 0],mem_1_0[0 + 1],mem_1_0[0 + 2],mem_1_0[0 + 3],mem_1_0[0 + 4],mem_1_0[0 + 5],mem_1_0[0 + 6],mem_1_0[0 + 7],mem_1_0[0 + 8],mem_1_0[0 + 9],mem_1_0[0 + 10],mem_1_0[0 + 11],mem_1_0[0 + 12],mem_1_0[0 + 13],mem_1_0[0 + 14],mem_1_0[0 + 15],mem_1_0[0 + 16],mem_1_0[0 + 17],mem_1_0[0 + 18],mem_1_0[0 + 19],mem_1_0[0 + 20],mem_1_0[0 + 21],mem_1_0[0 + 22],mem_1_0[0 + 23],mem_1_0[0 + 24],mem_1_0[0 + 25],mem_1_0[0 + 26],mem_1_0[0 + 27],mem_1_0[0 + 28],mem_1_0[0 + 29],mem_1_0[0 + 30],mem_1_0[0 + 31],mem_1_0[0 + 32],mem_1_0[0 + 33],mem_1_0[0 + 34],mem_1_0[0 + 35],mem_1_0[0 + 36],mem_1_0[0 + 37],mem_1_0[0 + 38],mem_1_0[0 + 39],mem_1_0[0 + 40],mem_1_0[0 + 41],mem_1_0[0 + 42],mem_1_0[0 + 43],mem_1_0[0 + 44],mem_1_0[0 + 45],mem_1_0[0 + 46],mem_1_0[0 + 47],mem_1_0[0 + 48],mem_1_0[0 + 49],mem_1_0[0 + 50],mem_1_0[0 + 51],mem_1_0[0 + 52],mem_1_0[0 + 53],mem_1_0[0 + 54],mem_1_0[0 + 55],mem_1_0[0 + 56],mem_1_0[0 + 57],mem_1_0[0 + 58],mem_1_0[0 + 59],mem_1_0[0 + 60],mem_1_0[0 + 61],mem_1_0[0 + 62],mem_1_0[0 + 63],mem_1_0[0 + 64],mem_1_0[0 + 65],mem_1_0[0 + 66],mem_1_0[0 + 67],mem_1_0[0 + 68],mem_1_0[0 + 69],mem_1_0[0 + 70],mem_1_0[0 + 71],mem_1_0[0 + 72],mem_1_0[0 + 73],mem_1_0[0 + 74],mem_1_0[0 + 75],mem_1_0[0 + 76],mem_1_0[0 + 77],mem_1_0[0 + 78],mem_1_0[0 + 79],mem_1_0[0 + 80],mem_1_0[0 + 81],mem_1_0[0 + 82],mem_1_0[0 + 83],mem_1_0[0 + 84],mem_1_0[0 + 85],mem_1_0[0 + 86],mem_1_0[0 + 87],mem_1_0[0 + 88],mem_1_0[0 + 89],mem_1_0[0 + 90],mem_1_0[0 + 91],mem_1_0[0 + 92],mem_1_0[0 + 93],mem_1_0[0 + 94],mem_1_0[0 + 95],mem_1_0[0 + 96],mem_1_0[0 + 97],mem_1_0[0 + 98],mem_1_0[0 + 99],mem_1_0[0 + 100],mem_1_0[0 + 101],mem_1_0[0 + 102],mem_1_0[0 + 103],mem_1_0[0 + 104],mem_1_0[0 + 105],mem_1_0[0 + 106],mem_1_0[0 + 107],mem_1_0[0 + 108],mem_1_0[0 + 109],mem_1_0[0 + 110],mem_1_0[0 + 111],mem_1_0[0 + 112],mem_1_0[0 + 113],mem_1_0[0 + 114],mem_1_0[0 + 115],mem_1_0[0 + 116],mem_1_0[0 + 117],mem_1_0[0 + 118],mem_1_0[0 + 119],mem_1_0[0 + 120],mem_1_0[0 + 121],mem_1_0[0 + 122],mem_1_0[0 + 123],mem_1_0[0 + 124],mem_1_0[0 + 125],mem_1_0[0 + 126],mem_1_0[0 + 127],mem_1_0[0 + 128],mem_1_0[0 + 129],mem_1_0[0 + 130],mem_1_0[0 + 131],mem_1_0[0 + 132],mem_1_0[0 + 133],mem_1_0[0 + 134],mem_1_0[0 + 135],mem_1_0[0 + 136],mem_1_0[0 + 137],mem_1_0[0 + 138],mem_1_0[0 + 139],mem_1_0[0 + 140],mem_1_0[0 + 141],mem_1_0[0 + 142],mem_1_0[0 + 143],mem_1_0[0 + 144],mem_1_0[0 + 145],mem_1_0[0 + 146],mem_1_0[0 + 147],mem_1_0[0 + 148],mem_1_0[0 + 149],mem_1_0[0 + 150],mem_1_0[0 + 151],mem_1_0[0 + 152],mem_1_0[0 + 153],mem_1_0[0 + 154],mem_1_0[0 + 155],mem_1_0[0 + 156],mem_1_0[0 + 157],mem_1_0[0 + 158],mem_1_0[0 + 159],mem_1_0[0 + 160],mem_1_0[0 + 161],mem_1_0[0 + 162],mem_1_0[0 + 163],mem_1_0[0 + 164],mem_1_0[0 + 165],mem_1_0[0 + 166],mem_1_0[0 + 167],mem_1_0[0 + 168],mem_1_0[0 + 169],mem_1_0[0 + 170],mem_1_0[0 + 171],mem_1_0[0 + 172],mem_1_0[0 + 173],mem_1_0[0 + 174],mem_1_0[0 + 175],mem_1_0[0 + 176],mem_1_0[0 + 177],mem_1_0[0 + 178],mem_1_0[0 + 179],mem_1_0[0 + 180],mem_1_0[0 + 181],mem_1_0[0 + 182],mem_1_0[0 + 183],mem_1_0[0 + 184],mem_1_0[0 + 185],mem_1_0[0 + 186],mem_1_0[0 + 187],mem_1_0[0 + 188],mem_1_0[0 + 189],mem_1_0[0 + 190],mem_1_0[0 + 191],mem_1_0[0 + 192],mem_1_0[0 + 193],mem_1_0[0 + 194],mem_1_0[0 + 195],mem_1_0[0 + 196],mem_1_0[0 + 197],mem_1_0[0 + 198],mem_1_0[0 + 199],mem_1_0[0 + 200],mem_1_0[0 + 201],mem_1_0[0 + 202],mem_1_0[0 + 203],mem_1_0[0 + 204],mem_1_0[0 + 205],mem_1_0[0 + 206],mem_1_0[0 + 207],mem_1_0[0 + 208],mem_1_0[0 + 209],mem_1_0[0 + 210],mem_1_0[0 + 211],mem_1_0[0 + 212],mem_1_0[0 + 213],mem_1_0[0 + 214],mem_1_0[0 + 215],mem_1_0[0 + 216],mem_1_0[0 + 217],mem_1_0[0 + 218],mem_1_0[0 + 219],mem_1_0[0 + 220],mem_1_0[0 + 221],mem_1_0[0 + 222],mem_1_0[0 + 223],mem_1_0[0 + 224],mem_1_0[0 + 225],mem_1_0[0 + 226],mem_1_0[0 + 227],mem_1_0[0 + 228],mem_1_0[0 + 229],mem_1_0[0 + 230],mem_1_0[0 + 231],mem_1_0[0 + 232],mem_1_0[0 + 233],mem_1_0[0 + 234],mem_1_0[0 + 235],mem_1_0[0 + 236],mem_1_0[0 + 237],mem_1_0[0 + 238],mem_1_0[0 + 239],mem_1_0[0 + 240],mem_1_0[0 + 241],mem_1_0[0 + 242],mem_1_0[0 + 243],mem_1_0[0 + 244],mem_1_0[0 + 245],mem_1_0[0 + 246],mem_1_0[0 + 247],mem_1_0[0 + 248],mem_1_0[0 + 249],mem_1_0[0 + 250],mem_1_0[0 + 251],mem_1_0[0 + 252],mem_1_0[0 + 253],mem_1_0[0 + 254],mem_1_0[0 + 255],mem_1_0[0 + 256],mem_1_0[0 + 257],mem_1_0[0 + 258],mem_1_0[0 + 259],mem_1_0[0 + 260],mem_1_0[0 + 261],mem_1_0[0 + 262],mem_1_0[0 + 263],mem_1_0[0 + 264],mem_1_0[0 + 265],mem_1_0[0 + 266],mem_1_0[0 + 267],mem_1_0[0 + 268],mem_1_0[0 + 269],mem_1_0[0 + 270],mem_1_0[0 + 271],mem_1_0[0 + 272],mem_1_0[0 + 273],mem_1_0[0 + 274],mem_1_0[0 + 275],mem_1_0[0 + 276],mem_1_0[0 + 277],mem_1_0[0 + 278],mem_1_0[0 + 279],mem_1_0[0 + 280],mem_1_0[0 + 281],mem_1_0[0 + 282],mem_1_0[0 + 283],mem_1_0[0 + 284],mem_1_0[0 + 285],mem_1_0[0 + 286],mem_1_0[0 + 287],mem_1_0[0 + 288],mem_1_0[0 + 289],mem_1_0[0 + 290],mem_1_0[0 + 291],mem_1_0[0 + 292],mem_1_0[0 + 293],mem_1_0[0 + 294],mem_1_0[0 + 295],mem_1_0[0 + 296],mem_1_0[0 + 297],mem_1_0[0 + 298],mem_1_0[0 + 299],mem_1_0[0 + 300],mem_1_0[0 + 301],mem_1_0[0 + 302],mem_1_0[0 + 303],mem_1_0[0 + 304],mem_1_0[0 + 305],mem_1_0[0 + 306],mem_1_0[0 + 307],mem_1_0[0 + 308],mem_1_0[0 + 309],mem_1_0[0 + 310],mem_1_0[0 + 311],mem_1_0[0 + 312],mem_1_0[0 + 313],mem_1_0[0 + 314],mem_1_0[0 + 315],mem_1_0[0 + 316],mem_1_0[0 + 317],mem_1_0[0 + 318],mem_1_0[0 + 319],mem_1_0[0 + 320],mem_1_0[0 + 321],mem_1_0[0 + 322],mem_1_0[0 + 323],mem_1_0[0 + 324],mem_1_0[0 + 325],mem_1_0[0 + 326],mem_1_0[0 + 327],mem_1_0[0 + 328],mem_1_0[0 + 329],mem_1_0[0 + 330],mem_1_0[0 + 331],mem_1_0[0 + 332],mem_1_0[0 + 333],mem_1_0[0 + 334],mem_1_0[0 + 335],mem_1_0[0 + 336],mem_1_0[0 + 337],mem_1_0[0 + 338],mem_1_0[0 + 339],mem_1_0[0 + 340],mem_1_0[0 + 341],mem_1_0[0 + 342],mem_1_0[0 + 343],mem_1_0[0 + 344],mem_1_0[0 + 345],mem_1_0[0 + 346],mem_1_0[0 + 347],mem_1_0[0 + 348],mem_1_0[0 + 349],mem_1_0[0 + 350],mem_1_0[0 + 351],mem_1_0[0 + 352],mem_1_0[0 + 353],mem_1_0[0 + 354],mem_1_0[0 + 355],mem_1_0[0 + 356],mem_1_0[0 + 357],mem_1_0[0 + 358],mem_1_0[0 + 359],mem_1_0[0 + 360],mem_1_0[0 + 361],mem_1_0[0 + 362],mem_1_0[0 + 363],mem_1_0[0 + 364],mem_1_0[0 + 365],mem_1_0[0 + 366],mem_1_0[0 + 367],mem_1_0[0 + 368],mem_1_0[0 + 369],mem_1_0[0 + 370],mem_1_0[0 + 371],mem_1_0[0 + 372],mem_1_0[0 + 373],mem_1_0[0 + 374],mem_1_0[0 + 375],mem_1_0[0 + 376],mem_1_0[0 + 377],mem_1_0[0 + 378],mem_1_0[0 + 379],mem_1_0[0 + 380],mem_1_0[0 + 381],mem_1_0[0 + 382],mem_1_0[0 + 383],mem_1_0[0 + 384],mem_1_0[0 + 385],mem_1_0[0 + 386],mem_1_0[0 + 387],mem_1_0[0 + 388],mem_1_0[0 + 389],mem_1_0[0 + 390],mem_1_0[0 + 391],mem_1_0[0 + 392],mem_1_0[0 + 393],mem_1_0[0 + 394],mem_1_0[0 + 395],mem_1_0[0 + 396],mem_1_0[0 + 397],mem_1_0[0 + 398],mem_1_0[0 + 399],mem_1_0[0 + 400],mem_1_0[0 + 401],mem_1_0[0 + 402],mem_1_0[0 + 403],mem_1_0[0 + 404],mem_1_0[0 + 405],mem_1_0[0 + 406],mem_1_0[0 + 407],mem_1_0[0 + 408],mem_1_0[0 + 409],mem_1_0[0 + 410],mem_1_0[0 + 411],mem_1_0[0 + 412],mem_1_0[0 + 413],mem_1_0[0 + 414],mem_1_0[0 + 415],mem_1_0[0 + 416],mem_1_0[0 + 417],mem_1_0[0 + 418],mem_1_0[0 + 419],mem_1_0[0 + 420],mem_1_0[0 + 421],mem_1_0[0 + 422],mem_1_0[0 + 423],mem_1_0[0 + 424],mem_1_0[0 + 425],mem_1_0[0 + 426],mem_1_0[0 + 427],mem_1_0[0 + 428],mem_1_0[0 + 429],mem_1_0[0 + 430],mem_1_0[0 + 431],mem_1_0[0 + 432],mem_1_0[0 + 433],mem_1_0[0 + 434],mem_1_0[0 + 435],mem_1_0[0 + 436],mem_1_0[0 + 437],mem_1_0[0 + 438],mem_1_0[0 + 439],mem_1_0[0 + 440],mem_1_0[0 + 441],mem_1_0[0 + 442],mem_1_0[0 + 443],mem_1_0[0 + 444],mem_1_0[0 + 445],mem_1_0[0 + 446],mem_1_0[0 + 447],mem_1_0[0 + 448],mem_1_0[0 + 449],mem_1_0[0 + 450],mem_1_0[0 + 451],mem_1_0[0 + 452],mem_1_0[0 + 453],mem_1_0[0 + 454],mem_1_0[0 + 455],mem_1_0[0 + 456],mem_1_0[0 + 457],mem_1_0[0 + 458],mem_1_0[0 + 459],mem_1_0[0 + 460],mem_1_0[0 + 461],mem_1_0[0 + 462],mem_1_0[0 + 463],mem_1_0[0 + 464],mem_1_0[0 + 465],mem_1_0[0 + 466],mem_1_0[0 + 467],mem_1_0[0 + 468],mem_1_0[0 + 469],mem_1_0[0 + 470],mem_1_0[0 + 471],mem_1_0[0 + 472],mem_1_0[0 + 473],mem_1_0[0 + 474],mem_1_0[0 + 475],mem_1_0[0 + 476],mem_1_0[0 + 477],mem_1_0[0 + 478],mem_1_0[0 + 479],mem_1_0[0 + 480],mem_1_0[0 + 481],mem_1_0[0 + 482],mem_1_0[0 + 483],mem_1_0[0 + 484],mem_1_0[0 + 485],mem_1_0[0 + 486],mem_1_0[0 + 487],mem_1_0[0 + 488],mem_1_0[0 + 489],mem_1_0[0 + 490],mem_1_0[0 + 491],mem_1_0[0 + 492],mem_1_0[0 + 493],mem_1_0[0 + 494],mem_1_0[0 + 495],mem_1_0[0 + 496],mem_1_0[0 + 497],mem_1_0[0 + 498],mem_1_0[0 + 499],mem_1_0[0 + 500],mem_1_0[0 + 501],mem_1_0[0 + 502],mem_1_0[0 + 503],mem_1_0[0 + 504],mem_1_0[0 + 505],mem_1_0[0 + 506],mem_1_0[0 + 507],mem_1_0[0 + 508],mem_1_0[0 + 509],mem_1_0[0 + 510],mem_1_0[0 + 511],mem_1_0[0 + 512],mem_1_0[0 + 513],mem_1_0[0 + 514],mem_1_0[0 + 515],mem_1_0[0 + 516],mem_1_0[0 + 517],mem_1_0[0 + 518],mem_1_0[0 + 519],mem_1_0[0 + 520],mem_1_0[0 + 521],mem_1_0[0 + 522],mem_1_0[0 + 523],mem_1_0[0 + 524],mem_1_0[0 + 525],mem_1_0[0 + 526],mem_1_0[0 + 527],mem_1_0[0 + 528],mem_1_0[0 + 529],mem_1_0[0 + 530],mem_1_0[0 + 531],mem_1_0[0 + 532],mem_1_0[0 + 533],mem_1_0[0 + 534],mem_1_0[0 + 535],mem_1_0[0 + 536],mem_1_0[0 + 537],mem_1_0[0 + 538],mem_1_0[0 + 539],mem_1_0[0 + 540],mem_1_0[0 + 541],mem_1_0[0 + 542],mem_1_0[0 + 543],mem_1_0[0 + 544],mem_1_0[0 + 545],mem_1_0[0 + 546],mem_1_0[0 + 547],mem_1_0[0 + 548],mem_1_0[0 + 549],mem_1_0[0 + 550],mem_1_0[0 + 551],mem_1_0[0 + 552],mem_1_0[0 + 553],mem_1_0[0 + 554],mem_1_0[0 + 555],mem_1_0[0 + 556],mem_1_0[0 + 557],mem_1_0[0 + 558],mem_1_0[0 + 559],mem_1_0[0 + 560],mem_1_0[0 + 561],mem_1_0[0 + 562],mem_1_0[0 + 563],mem_1_0[0 + 564],mem_1_0[0 + 565],mem_1_0[0 + 566],mem_1_0[0 + 567],mem_1_0[0 + 568],mem_1_0[0 + 569],mem_1_0[0 + 570],mem_1_0[0 + 571],mem_1_0[0 + 572],mem_1_0[0 + 573],mem_1_0[0 + 574],mem_1_0[0 + 575],mem_1_0[0 + 576],mem_1_0[0 + 577],mem_1_0[0 + 578],mem_1_0[0 + 579],mem_1_0[0 + 580],mem_1_0[0 + 581],mem_1_0[0 + 582],mem_1_0[0 + 583],mem_1_0[0 + 584],mem_1_0[0 + 585],mem_1_0[0 + 586],mem_1_0[0 + 587],mem_1_0[0 + 588],mem_1_0[0 + 589],mem_1_0[0 + 590],mem_1_0[0 + 591],mem_1_0[0 + 592],mem_1_0[0 + 593],mem_1_0[0 + 594],mem_1_0[0 + 595],mem_1_0[0 + 596],mem_1_0[0 + 597],mem_1_0[0 + 598],mem_1_0[0 + 599],mem_1_0[0 + 600],mem_1_0[0 + 601],mem_1_0[0 + 602],mem_1_0[0 + 603],mem_1_0[0 + 604],mem_1_0[0 + 605],mem_1_0[0 + 606],mem_1_0[0 + 607],mem_1_0[0 + 608],mem_1_0[0 + 609],mem_1_0[0 + 610],mem_1_0[0 + 611],mem_1_0[0 + 612],mem_1_0[0 + 613],mem_1_0[0 + 614],mem_1_0[0 + 615],mem_1_0[0 + 616],mem_1_0[0 + 617],mem_1_0[0 + 618],mem_1_0[0 + 619],mem_1_0[0 + 620],mem_1_0[0 + 621],mem_1_0[0 + 622],mem_1_0[0 + 623],mem_1_0[0 + 624],mem_1_0[0 + 625],mem_1_0[0 + 626],mem_1_0[0 + 627],mem_1_0[0 + 628],mem_1_0[0 + 629],mem_1_0[0 + 630],mem_1_0[0 + 631],mem_1_0[0 + 632],mem_1_0[0 + 633],mem_1_0[0 + 634],mem_1_0[0 + 635],mem_1_0[0 + 636],mem_1_0[0 + 637],mem_1_0[0 + 638],mem_1_0[0 + 639],mem_1_0[0 + 640],mem_1_0[0 + 641],mem_1_0[0 + 642],mem_1_0[0 + 643],mem_1_0[0 + 644],mem_1_0[0 + 645],mem_1_0[0 + 646],mem_1_0[0 + 647],mem_1_0[0 + 648],mem_1_0[0 + 649],mem_1_0[0 + 650],mem_1_0[0 + 651],mem_1_0[0 + 652],mem_1_0[0 + 653],mem_1_0[0 + 654],mem_1_0[0 + 655],mem_1_0[0 + 656],mem_1_0[0 + 657],mem_1_0[0 + 658],mem_1_0[0 + 659],mem_1_0[0 + 660],mem_1_0[0 + 661],mem_1_0[0 + 662],mem_1_0[0 + 663],mem_1_0[0 + 664],mem_1_0[0 + 665],mem_1_0[0 + 666],mem_1_0[0 + 667],mem_1_0[0 + 668],mem_1_0[0 + 669],mem_1_0[0 + 670],mem_1_0[0 + 671],mem_1_0[0 + 672],mem_1_0[0 + 673],mem_1_0[0 + 674],mem_1_0[0 + 675],mem_1_0[0 + 676],mem_1_0[0 + 677],mem_1_0[0 + 678],mem_1_0[0 + 679],mem_1_0[0 + 680],mem_1_0[0 + 681],mem_1_0[0 + 682],mem_1_0[0 + 683],mem_1_0[0 + 684],mem_1_0[0 + 685],mem_1_0[0 + 686],mem_1_0[0 + 687],mem_1_0[0 + 688],mem_1_0[0 + 689],mem_1_0[0 + 690],mem_1_0[0 + 691],mem_1_0[0 + 692],mem_1_0[0 + 693],mem_1_0[0 + 694],mem_1_0[0 + 695],mem_1_0[0 + 696],mem_1_0[0 + 697],mem_1_0[0 + 698],mem_1_0[0 + 699],mem_1_0[0 + 700],mem_1_0[0 + 701],mem_1_0[0 + 702],mem_1_0[0 + 703],mem_1_0[0 + 704],mem_1_0[0 + 705],mem_1_0[0 + 706],mem_1_0[0 + 707],mem_1_0[0 + 708],mem_1_0[0 + 709],mem_1_0[0 + 710],mem_1_0[0 + 711],mem_1_0[0 + 712],mem_1_0[0 + 713],mem_1_0[0 + 714],mem_1_0[0 + 715],mem_1_0[0 + 716],mem_1_0[0 + 717],mem_1_0[0 + 718],mem_1_0[0 + 719],mem_1_0[0 + 720],mem_1_0[0 + 721],mem_1_0[0 + 722],mem_1_0[0 + 723],mem_1_0[0 + 724],mem_1_0[0 + 725],mem_1_0[0 + 726],mem_1_0[0 + 727],mem_1_0[0 + 728],mem_1_0[0 + 729],mem_1_0[0 + 730],mem_1_0[0 + 731],mem_1_0[0 + 732],mem_1_0[0 + 733],mem_1_0[0 + 734],mem_1_0[0 + 735],mem_1_0[0 + 736],mem_1_0[0 + 737],mem_1_0[0 + 738],mem_1_0[0 + 739],mem_1_0[0 + 740],mem_1_0[0 + 741],mem_1_0[0 + 742],mem_1_0[0 + 743],mem_1_0[0 + 744],mem_1_0[0 + 745],mem_1_0[0 + 746],mem_1_0[0 + 747],mem_1_0[0 + 748],mem_1_0[0 + 749],mem_1_0[0 + 750],mem_1_0[0 + 751],mem_1_0[0 + 752],mem_1_0[0 + 753],mem_1_0[0 + 754],mem_1_0[0 + 755],mem_1_0[0 + 756],mem_1_0[0 + 757],mem_1_0[0 + 758],mem_1_0[0 + 759],mem_1_0[0 + 760],mem_1_0[0 + 761],mem_1_0[0 + 762],mem_1_0[0 + 763],mem_1_0[0 + 764],mem_1_0[0 + 765],mem_1_0[0 + 766],mem_1_0[0 + 767],mem_1_0[0 + 768],mem_1_0[0 + 769],mem_1_0[0 + 770],mem_1_0[0 + 771],mem_1_0[0 + 772],mem_1_0[0 + 773],mem_1_0[0 + 774],mem_1_0[0 + 775],mem_1_0[0 + 776],mem_1_0[0 + 777],mem_1_0[0 + 778],mem_1_0[0 + 779],mem_1_0[0 + 780],mem_1_0[0 + 781],mem_1_0[0 + 782],mem_1_0[0 + 783],mem_1_0[0 + 784],mem_1_0[0 + 785],mem_1_0[0 + 786],mem_1_0[0 + 787],mem_1_0[0 + 788],mem_1_0[0 + 789],mem_1_0[0 + 790],mem_1_0[0 + 791],mem_1_0[0 + 792],mem_1_0[0 + 793],mem_1_0[0 + 794],mem_1_0[0 + 795],mem_1_0[0 + 796],mem_1_0[0 + 797],mem_1_0[0 + 798],mem_1_0[0 + 799],mem_1_0[0 + 800],mem_1_0[0 + 801],mem_1_0[0 + 802],mem_1_0[0 + 803],mem_1_0[0 + 804],mem_1_0[0 + 805],mem_1_0[0 + 806],mem_1_0[0 + 807],mem_1_0[0 + 808],mem_1_0[0 + 809],mem_1_0[0 + 810],mem_1_0[0 + 811],mem_1_0[0 + 812],mem_1_0[0 + 813],mem_1_0[0 + 814],mem_1_0[0 + 815],mem_1_0[0 + 816],mem_1_0[0 + 817],mem_1_0[0 + 818],mem_1_0[0 + 819],mem_1_0[0 + 820],mem_1_0[0 + 821],mem_1_0[0 + 822],mem_1_0[0 + 823],mem_1_0[0 + 824],mem_1_0[0 + 825],mem_1_0[0 + 826],mem_1_0[0 + 827],mem_1_0[0 + 828],mem_1_0[0 + 829],mem_1_0[0 + 830],mem_1_0[0 + 831],mem_1_0[0 + 832],mem_1_0[0 + 833],mem_1_0[0 + 834],mem_1_0[0 + 835],mem_1_0[0 + 836],mem_1_0[0 + 837],mem_1_0[0 + 838],mem_1_0[0 + 839],mem_1_0[0 + 840],mem_1_0[0 + 841],mem_1_0[0 + 842],mem_1_0[0 + 843],mem_1_0[0 + 844],mem_1_0[0 + 845],mem_1_0[0 + 846],mem_1_0[0 + 847],mem_1_0[0 + 848],mem_1_0[0 + 849],mem_1_0[0 + 850],mem_1_0[0 + 851],mem_1_0[0 + 852],mem_1_0[0 + 853],mem_1_0[0 + 854],mem_1_0[0 + 855],mem_1_0[0 + 856],mem_1_0[0 + 857],mem_1_0[0 + 858],mem_1_0[0 + 859],mem_1_0[0 + 860],mem_1_0[0 + 861],mem_1_0[0 + 862],mem_1_0[0 + 863],mem_1_0[0 + 864],mem_1_0[0 + 865],mem_1_0[0 + 866],mem_1_0[0 + 867],mem_1_0[0 + 868],mem_1_0[0 + 869],mem_1_0[0 + 870],mem_1_0[0 + 871],mem_1_0[0 + 872],mem_1_0[0 + 873],mem_1_0[0 + 874],mem_1_0[0 + 875],mem_1_0[0 + 876],mem_1_0[0 + 877],mem_1_0[0 + 878],mem_1_0[0 + 879],mem_1_0[0 + 880],mem_1_0[0 + 881],mem_1_0[0 + 882],mem_1_0[0 + 883],mem_1_0[0 + 884],mem_1_0[0 + 885],mem_1_0[0 + 886],mem_1_0[0 + 887],mem_1_0[0 + 888],mem_1_0[0 + 889],mem_1_0[0 + 890],mem_1_0[0 + 891],mem_1_0[0 + 892],mem_1_0[0 + 893],mem_1_0[0 + 894],mem_1_0[0 + 895],mem_1_0[0 + 896],mem_1_0[0 + 897],mem_1_0[0 + 898],mem_1_0[0 + 899],mem_1_0[0 + 900],mem_1_0[0 + 901],mem_1_0[0 + 902],mem_1_0[0 + 903],mem_1_0[0 + 904],mem_1_0[0 + 905],mem_1_0[0 + 906],mem_1_0[0 + 907],mem_1_0[0 + 908],mem_1_0[0 + 909],mem_1_0[0 + 910],mem_1_0[0 + 911],mem_1_0[0 + 912],mem_1_0[0 + 913],mem_1_0[0 + 914],mem_1_0[0 + 915],mem_1_0[0 + 916],mem_1_0[0 + 917],mem_1_0[0 + 918],mem_1_0[0 + 919],mem_1_0[0 + 920],mem_1_0[0 + 921],mem_1_0[0 + 922],mem_1_0[0 + 923],mem_1_0[0 + 924],mem_1_0[0 + 925],mem_1_0[0 + 926],mem_1_0[0 + 927],mem_1_0[0 + 928],mem_1_0[0 + 929],mem_1_0[0 + 930],mem_1_0[0 + 931],mem_1_0[0 + 932],mem_1_0[0 + 933],mem_1_0[0 + 934],mem_1_0[0 + 935],mem_1_0[0 + 936],mem_1_0[0 + 937],mem_1_0[0 + 938],mem_1_0[0 + 939],mem_1_0[0 + 940],mem_1_0[0 + 941],mem_1_0[0 + 942],mem_1_0[0 + 943],mem_1_0[0 + 944],mem_1_0[0 + 945],mem_1_0[0 + 946],mem_1_0[0 + 947],mem_1_0[0 + 948],mem_1_0[0 + 949],mem_1_0[0 + 950],mem_1_0[0 + 951],mem_1_0[0 + 952],mem_1_0[0 + 953],mem_1_0[0 + 954],mem_1_0[0 + 955],mem_1_0[0 + 956],mem_1_0[0 + 957],mem_1_0[0 + 958],mem_1_0[0 + 959],mem_1_0[0 + 960],mem_1_0[0 + 961],mem_1_0[0 + 962],mem_1_0[0 + 963],mem_1_0[0 + 964],mem_1_0[0 + 965],mem_1_0[0 + 966],mem_1_0[0 + 967],mem_1_0[0 + 968],mem_1_0[0 + 969],mem_1_0[0 + 970],mem_1_0[0 + 971],mem_1_0[0 + 972],mem_1_0[0 + 973],mem_1_0[0 + 974],mem_1_0[0 + 975],mem_1_0[0 + 976],mem_1_0[0 + 977],mem_1_0[0 + 978],mem_1_0[0 + 979],mem_1_0[0 + 980],mem_1_0[0 + 981],mem_1_0[0 + 982],mem_1_0[0 + 983],mem_1_0[0 + 984],mem_1_0[0 + 985],mem_1_0[0 + 986],mem_1_0[0 + 987],mem_1_0[0 + 988],mem_1_0[0 + 989],mem_1_0[0 + 990],mem_1_0[0 + 991],mem_1_0[0 + 992],mem_1_0[0 + 993],mem_1_0[0 + 994],mem_1_0[0 + 995],mem_1_0[0 + 996],mem_1_0[0 + 997],mem_1_0[0 + 998],mem_1_0[0 + 999],mem_1_0[0 + 1000],mem_1_0[0 + 1001],mem_1_0[0 + 1002],mem_1_0[0 + 1003],mem_1_0[0 + 1004],mem_1_0[0 + 1005],mem_1_0[0 + 1006],mem_1_0[0 + 1007],mem_1_0[0 + 1008],mem_1_0[0 + 1009],mem_1_0[0 + 1010],mem_1_0[0 + 1011],mem_1_0[0 + 1012],mem_1_0[0 + 1013],mem_1_0[0 + 1014],mem_1_0[0 + 1015],mem_1_0[0 + 1016],mem_1_0[0 + 1017],mem_1_0[0 + 1018],mem_1_0[0 + 1019],mem_1_0[0 + 1020],mem_1_0[0 + 1021],mem_1_0[0 + 1022],mem_1_0[0 + 1024 - 1] };
wire [8*(1024)-1:0] mem_2_0_flat_src;
assign mem_2_0_flat_src = {mem_2_0[0 + 0],mem_2_0[0 + 1],mem_2_0[0 + 2],mem_2_0[0 + 3],mem_2_0[0 + 4],mem_2_0[0 + 5],mem_2_0[0 + 6],mem_2_0[0 + 7],mem_2_0[0 + 8],mem_2_0[0 + 9],mem_2_0[0 + 10],mem_2_0[0 + 11],mem_2_0[0 + 12],mem_2_0[0 + 13],mem_2_0[0 + 14],mem_2_0[0 + 15],mem_2_0[0 + 16],mem_2_0[0 + 17],mem_2_0[0 + 18],mem_2_0[0 + 19],mem_2_0[0 + 20],mem_2_0[0 + 21],mem_2_0[0 + 22],mem_2_0[0 + 23],mem_2_0[0 + 24],mem_2_0[0 + 25],mem_2_0[0 + 26],mem_2_0[0 + 27],mem_2_0[0 + 28],mem_2_0[0 + 29],mem_2_0[0 + 30],mem_2_0[0 + 31],mem_2_0[0 + 32],mem_2_0[0 + 33],mem_2_0[0 + 34],mem_2_0[0 + 35],mem_2_0[0 + 36],mem_2_0[0 + 37],mem_2_0[0 + 38],mem_2_0[0 + 39],mem_2_0[0 + 40],mem_2_0[0 + 41],mem_2_0[0 + 42],mem_2_0[0 + 43],mem_2_0[0 + 44],mem_2_0[0 + 45],mem_2_0[0 + 46],mem_2_0[0 + 47],mem_2_0[0 + 48],mem_2_0[0 + 49],mem_2_0[0 + 50],mem_2_0[0 + 51],mem_2_0[0 + 52],mem_2_0[0 + 53],mem_2_0[0 + 54],mem_2_0[0 + 55],mem_2_0[0 + 56],mem_2_0[0 + 57],mem_2_0[0 + 58],mem_2_0[0 + 59],mem_2_0[0 + 60],mem_2_0[0 + 61],mem_2_0[0 + 62],mem_2_0[0 + 63],mem_2_0[0 + 64],mem_2_0[0 + 65],mem_2_0[0 + 66],mem_2_0[0 + 67],mem_2_0[0 + 68],mem_2_0[0 + 69],mem_2_0[0 + 70],mem_2_0[0 + 71],mem_2_0[0 + 72],mem_2_0[0 + 73],mem_2_0[0 + 74],mem_2_0[0 + 75],mem_2_0[0 + 76],mem_2_0[0 + 77],mem_2_0[0 + 78],mem_2_0[0 + 79],mem_2_0[0 + 80],mem_2_0[0 + 81],mem_2_0[0 + 82],mem_2_0[0 + 83],mem_2_0[0 + 84],mem_2_0[0 + 85],mem_2_0[0 + 86],mem_2_0[0 + 87],mem_2_0[0 + 88],mem_2_0[0 + 89],mem_2_0[0 + 90],mem_2_0[0 + 91],mem_2_0[0 + 92],mem_2_0[0 + 93],mem_2_0[0 + 94],mem_2_0[0 + 95],mem_2_0[0 + 96],mem_2_0[0 + 97],mem_2_0[0 + 98],mem_2_0[0 + 99],mem_2_0[0 + 100],mem_2_0[0 + 101],mem_2_0[0 + 102],mem_2_0[0 + 103],mem_2_0[0 + 104],mem_2_0[0 + 105],mem_2_0[0 + 106],mem_2_0[0 + 107],mem_2_0[0 + 108],mem_2_0[0 + 109],mem_2_0[0 + 110],mem_2_0[0 + 111],mem_2_0[0 + 112],mem_2_0[0 + 113],mem_2_0[0 + 114],mem_2_0[0 + 115],mem_2_0[0 + 116],mem_2_0[0 + 117],mem_2_0[0 + 118],mem_2_0[0 + 119],mem_2_0[0 + 120],mem_2_0[0 + 121],mem_2_0[0 + 122],mem_2_0[0 + 123],mem_2_0[0 + 124],mem_2_0[0 + 125],mem_2_0[0 + 126],mem_2_0[0 + 127],mem_2_0[0 + 128],mem_2_0[0 + 129],mem_2_0[0 + 130],mem_2_0[0 + 131],mem_2_0[0 + 132],mem_2_0[0 + 133],mem_2_0[0 + 134],mem_2_0[0 + 135],mem_2_0[0 + 136],mem_2_0[0 + 137],mem_2_0[0 + 138],mem_2_0[0 + 139],mem_2_0[0 + 140],mem_2_0[0 + 141],mem_2_0[0 + 142],mem_2_0[0 + 143],mem_2_0[0 + 144],mem_2_0[0 + 145],mem_2_0[0 + 146],mem_2_0[0 + 147],mem_2_0[0 + 148],mem_2_0[0 + 149],mem_2_0[0 + 150],mem_2_0[0 + 151],mem_2_0[0 + 152],mem_2_0[0 + 153],mem_2_0[0 + 154],mem_2_0[0 + 155],mem_2_0[0 + 156],mem_2_0[0 + 157],mem_2_0[0 + 158],mem_2_0[0 + 159],mem_2_0[0 + 160],mem_2_0[0 + 161],mem_2_0[0 + 162],mem_2_0[0 + 163],mem_2_0[0 + 164],mem_2_0[0 + 165],mem_2_0[0 + 166],mem_2_0[0 + 167],mem_2_0[0 + 168],mem_2_0[0 + 169],mem_2_0[0 + 170],mem_2_0[0 + 171],mem_2_0[0 + 172],mem_2_0[0 + 173],mem_2_0[0 + 174],mem_2_0[0 + 175],mem_2_0[0 + 176],mem_2_0[0 + 177],mem_2_0[0 + 178],mem_2_0[0 + 179],mem_2_0[0 + 180],mem_2_0[0 + 181],mem_2_0[0 + 182],mem_2_0[0 + 183],mem_2_0[0 + 184],mem_2_0[0 + 185],mem_2_0[0 + 186],mem_2_0[0 + 187],mem_2_0[0 + 188],mem_2_0[0 + 189],mem_2_0[0 + 190],mem_2_0[0 + 191],mem_2_0[0 + 192],mem_2_0[0 + 193],mem_2_0[0 + 194],mem_2_0[0 + 195],mem_2_0[0 + 196],mem_2_0[0 + 197],mem_2_0[0 + 198],mem_2_0[0 + 199],mem_2_0[0 + 200],mem_2_0[0 + 201],mem_2_0[0 + 202],mem_2_0[0 + 203],mem_2_0[0 + 204],mem_2_0[0 + 205],mem_2_0[0 + 206],mem_2_0[0 + 207],mem_2_0[0 + 208],mem_2_0[0 + 209],mem_2_0[0 + 210],mem_2_0[0 + 211],mem_2_0[0 + 212],mem_2_0[0 + 213],mem_2_0[0 + 214],mem_2_0[0 + 215],mem_2_0[0 + 216],mem_2_0[0 + 217],mem_2_0[0 + 218],mem_2_0[0 + 219],mem_2_0[0 + 220],mem_2_0[0 + 221],mem_2_0[0 + 222],mem_2_0[0 + 223],mem_2_0[0 + 224],mem_2_0[0 + 225],mem_2_0[0 + 226],mem_2_0[0 + 227],mem_2_0[0 + 228],mem_2_0[0 + 229],mem_2_0[0 + 230],mem_2_0[0 + 231],mem_2_0[0 + 232],mem_2_0[0 + 233],mem_2_0[0 + 234],mem_2_0[0 + 235],mem_2_0[0 + 236],mem_2_0[0 + 237],mem_2_0[0 + 238],mem_2_0[0 + 239],mem_2_0[0 + 240],mem_2_0[0 + 241],mem_2_0[0 + 242],mem_2_0[0 + 243],mem_2_0[0 + 244],mem_2_0[0 + 245],mem_2_0[0 + 246],mem_2_0[0 + 247],mem_2_0[0 + 248],mem_2_0[0 + 249],mem_2_0[0 + 250],mem_2_0[0 + 251],mem_2_0[0 + 252],mem_2_0[0 + 253],mem_2_0[0 + 254],mem_2_0[0 + 255],mem_2_0[0 + 256],mem_2_0[0 + 257],mem_2_0[0 + 258],mem_2_0[0 + 259],mem_2_0[0 + 260],mem_2_0[0 + 261],mem_2_0[0 + 262],mem_2_0[0 + 263],mem_2_0[0 + 264],mem_2_0[0 + 265],mem_2_0[0 + 266],mem_2_0[0 + 267],mem_2_0[0 + 268],mem_2_0[0 + 269],mem_2_0[0 + 270],mem_2_0[0 + 271],mem_2_0[0 + 272],mem_2_0[0 + 273],mem_2_0[0 + 274],mem_2_0[0 + 275],mem_2_0[0 + 276],mem_2_0[0 + 277],mem_2_0[0 + 278],mem_2_0[0 + 279],mem_2_0[0 + 280],mem_2_0[0 + 281],mem_2_0[0 + 282],mem_2_0[0 + 283],mem_2_0[0 + 284],mem_2_0[0 + 285],mem_2_0[0 + 286],mem_2_0[0 + 287],mem_2_0[0 + 288],mem_2_0[0 + 289],mem_2_0[0 + 290],mem_2_0[0 + 291],mem_2_0[0 + 292],mem_2_0[0 + 293],mem_2_0[0 + 294],mem_2_0[0 + 295],mem_2_0[0 + 296],mem_2_0[0 + 297],mem_2_0[0 + 298],mem_2_0[0 + 299],mem_2_0[0 + 300],mem_2_0[0 + 301],mem_2_0[0 + 302],mem_2_0[0 + 303],mem_2_0[0 + 304],mem_2_0[0 + 305],mem_2_0[0 + 306],mem_2_0[0 + 307],mem_2_0[0 + 308],mem_2_0[0 + 309],mem_2_0[0 + 310],mem_2_0[0 + 311],mem_2_0[0 + 312],mem_2_0[0 + 313],mem_2_0[0 + 314],mem_2_0[0 + 315],mem_2_0[0 + 316],mem_2_0[0 + 317],mem_2_0[0 + 318],mem_2_0[0 + 319],mem_2_0[0 + 320],mem_2_0[0 + 321],mem_2_0[0 + 322],mem_2_0[0 + 323],mem_2_0[0 + 324],mem_2_0[0 + 325],mem_2_0[0 + 326],mem_2_0[0 + 327],mem_2_0[0 + 328],mem_2_0[0 + 329],mem_2_0[0 + 330],mem_2_0[0 + 331],mem_2_0[0 + 332],mem_2_0[0 + 333],mem_2_0[0 + 334],mem_2_0[0 + 335],mem_2_0[0 + 336],mem_2_0[0 + 337],mem_2_0[0 + 338],mem_2_0[0 + 339],mem_2_0[0 + 340],mem_2_0[0 + 341],mem_2_0[0 + 342],mem_2_0[0 + 343],mem_2_0[0 + 344],mem_2_0[0 + 345],mem_2_0[0 + 346],mem_2_0[0 + 347],mem_2_0[0 + 348],mem_2_0[0 + 349],mem_2_0[0 + 350],mem_2_0[0 + 351],mem_2_0[0 + 352],mem_2_0[0 + 353],mem_2_0[0 + 354],mem_2_0[0 + 355],mem_2_0[0 + 356],mem_2_0[0 + 357],mem_2_0[0 + 358],mem_2_0[0 + 359],mem_2_0[0 + 360],mem_2_0[0 + 361],mem_2_0[0 + 362],mem_2_0[0 + 363],mem_2_0[0 + 364],mem_2_0[0 + 365],mem_2_0[0 + 366],mem_2_0[0 + 367],mem_2_0[0 + 368],mem_2_0[0 + 369],mem_2_0[0 + 370],mem_2_0[0 + 371],mem_2_0[0 + 372],mem_2_0[0 + 373],mem_2_0[0 + 374],mem_2_0[0 + 375],mem_2_0[0 + 376],mem_2_0[0 + 377],mem_2_0[0 + 378],mem_2_0[0 + 379],mem_2_0[0 + 380],mem_2_0[0 + 381],mem_2_0[0 + 382],mem_2_0[0 + 383],mem_2_0[0 + 384],mem_2_0[0 + 385],mem_2_0[0 + 386],mem_2_0[0 + 387],mem_2_0[0 + 388],mem_2_0[0 + 389],mem_2_0[0 + 390],mem_2_0[0 + 391],mem_2_0[0 + 392],mem_2_0[0 + 393],mem_2_0[0 + 394],mem_2_0[0 + 395],mem_2_0[0 + 396],mem_2_0[0 + 397],mem_2_0[0 + 398],mem_2_0[0 + 399],mem_2_0[0 + 400],mem_2_0[0 + 401],mem_2_0[0 + 402],mem_2_0[0 + 403],mem_2_0[0 + 404],mem_2_0[0 + 405],mem_2_0[0 + 406],mem_2_0[0 + 407],mem_2_0[0 + 408],mem_2_0[0 + 409],mem_2_0[0 + 410],mem_2_0[0 + 411],mem_2_0[0 + 412],mem_2_0[0 + 413],mem_2_0[0 + 414],mem_2_0[0 + 415],mem_2_0[0 + 416],mem_2_0[0 + 417],mem_2_0[0 + 418],mem_2_0[0 + 419],mem_2_0[0 + 420],mem_2_0[0 + 421],mem_2_0[0 + 422],mem_2_0[0 + 423],mem_2_0[0 + 424],mem_2_0[0 + 425],mem_2_0[0 + 426],mem_2_0[0 + 427],mem_2_0[0 + 428],mem_2_0[0 + 429],mem_2_0[0 + 430],mem_2_0[0 + 431],mem_2_0[0 + 432],mem_2_0[0 + 433],mem_2_0[0 + 434],mem_2_0[0 + 435],mem_2_0[0 + 436],mem_2_0[0 + 437],mem_2_0[0 + 438],mem_2_0[0 + 439],mem_2_0[0 + 440],mem_2_0[0 + 441],mem_2_0[0 + 442],mem_2_0[0 + 443],mem_2_0[0 + 444],mem_2_0[0 + 445],mem_2_0[0 + 446],mem_2_0[0 + 447],mem_2_0[0 + 448],mem_2_0[0 + 449],mem_2_0[0 + 450],mem_2_0[0 + 451],mem_2_0[0 + 452],mem_2_0[0 + 453],mem_2_0[0 + 454],mem_2_0[0 + 455],mem_2_0[0 + 456],mem_2_0[0 + 457],mem_2_0[0 + 458],mem_2_0[0 + 459],mem_2_0[0 + 460],mem_2_0[0 + 461],mem_2_0[0 + 462],mem_2_0[0 + 463],mem_2_0[0 + 464],mem_2_0[0 + 465],mem_2_0[0 + 466],mem_2_0[0 + 467],mem_2_0[0 + 468],mem_2_0[0 + 469],mem_2_0[0 + 470],mem_2_0[0 + 471],mem_2_0[0 + 472],mem_2_0[0 + 473],mem_2_0[0 + 474],mem_2_0[0 + 475],mem_2_0[0 + 476],mem_2_0[0 + 477],mem_2_0[0 + 478],mem_2_0[0 + 479],mem_2_0[0 + 480],mem_2_0[0 + 481],mem_2_0[0 + 482],mem_2_0[0 + 483],mem_2_0[0 + 484],mem_2_0[0 + 485],mem_2_0[0 + 486],mem_2_0[0 + 487],mem_2_0[0 + 488],mem_2_0[0 + 489],mem_2_0[0 + 490],mem_2_0[0 + 491],mem_2_0[0 + 492],mem_2_0[0 + 493],mem_2_0[0 + 494],mem_2_0[0 + 495],mem_2_0[0 + 496],mem_2_0[0 + 497],mem_2_0[0 + 498],mem_2_0[0 + 499],mem_2_0[0 + 500],mem_2_0[0 + 501],mem_2_0[0 + 502],mem_2_0[0 + 503],mem_2_0[0 + 504],mem_2_0[0 + 505],mem_2_0[0 + 506],mem_2_0[0 + 507],mem_2_0[0 + 508],mem_2_0[0 + 509],mem_2_0[0 + 510],mem_2_0[0 + 511],mem_2_0[0 + 512],mem_2_0[0 + 513],mem_2_0[0 + 514],mem_2_0[0 + 515],mem_2_0[0 + 516],mem_2_0[0 + 517],mem_2_0[0 + 518],mem_2_0[0 + 519],mem_2_0[0 + 520],mem_2_0[0 + 521],mem_2_0[0 + 522],mem_2_0[0 + 523],mem_2_0[0 + 524],mem_2_0[0 + 525],mem_2_0[0 + 526],mem_2_0[0 + 527],mem_2_0[0 + 528],mem_2_0[0 + 529],mem_2_0[0 + 530],mem_2_0[0 + 531],mem_2_0[0 + 532],mem_2_0[0 + 533],mem_2_0[0 + 534],mem_2_0[0 + 535],mem_2_0[0 + 536],mem_2_0[0 + 537],mem_2_0[0 + 538],mem_2_0[0 + 539],mem_2_0[0 + 540],mem_2_0[0 + 541],mem_2_0[0 + 542],mem_2_0[0 + 543],mem_2_0[0 + 544],mem_2_0[0 + 545],mem_2_0[0 + 546],mem_2_0[0 + 547],mem_2_0[0 + 548],mem_2_0[0 + 549],mem_2_0[0 + 550],mem_2_0[0 + 551],mem_2_0[0 + 552],mem_2_0[0 + 553],mem_2_0[0 + 554],mem_2_0[0 + 555],mem_2_0[0 + 556],mem_2_0[0 + 557],mem_2_0[0 + 558],mem_2_0[0 + 559],mem_2_0[0 + 560],mem_2_0[0 + 561],mem_2_0[0 + 562],mem_2_0[0 + 563],mem_2_0[0 + 564],mem_2_0[0 + 565],mem_2_0[0 + 566],mem_2_0[0 + 567],mem_2_0[0 + 568],mem_2_0[0 + 569],mem_2_0[0 + 570],mem_2_0[0 + 571],mem_2_0[0 + 572],mem_2_0[0 + 573],mem_2_0[0 + 574],mem_2_0[0 + 575],mem_2_0[0 + 576],mem_2_0[0 + 577],mem_2_0[0 + 578],mem_2_0[0 + 579],mem_2_0[0 + 580],mem_2_0[0 + 581],mem_2_0[0 + 582],mem_2_0[0 + 583],mem_2_0[0 + 584],mem_2_0[0 + 585],mem_2_0[0 + 586],mem_2_0[0 + 587],mem_2_0[0 + 588],mem_2_0[0 + 589],mem_2_0[0 + 590],mem_2_0[0 + 591],mem_2_0[0 + 592],mem_2_0[0 + 593],mem_2_0[0 + 594],mem_2_0[0 + 595],mem_2_0[0 + 596],mem_2_0[0 + 597],mem_2_0[0 + 598],mem_2_0[0 + 599],mem_2_0[0 + 600],mem_2_0[0 + 601],mem_2_0[0 + 602],mem_2_0[0 + 603],mem_2_0[0 + 604],mem_2_0[0 + 605],mem_2_0[0 + 606],mem_2_0[0 + 607],mem_2_0[0 + 608],mem_2_0[0 + 609],mem_2_0[0 + 610],mem_2_0[0 + 611],mem_2_0[0 + 612],mem_2_0[0 + 613],mem_2_0[0 + 614],mem_2_0[0 + 615],mem_2_0[0 + 616],mem_2_0[0 + 617],mem_2_0[0 + 618],mem_2_0[0 + 619],mem_2_0[0 + 620],mem_2_0[0 + 621],mem_2_0[0 + 622],mem_2_0[0 + 623],mem_2_0[0 + 624],mem_2_0[0 + 625],mem_2_0[0 + 626],mem_2_0[0 + 627],mem_2_0[0 + 628],mem_2_0[0 + 629],mem_2_0[0 + 630],mem_2_0[0 + 631],mem_2_0[0 + 632],mem_2_0[0 + 633],mem_2_0[0 + 634],mem_2_0[0 + 635],mem_2_0[0 + 636],mem_2_0[0 + 637],mem_2_0[0 + 638],mem_2_0[0 + 639],mem_2_0[0 + 640],mem_2_0[0 + 641],mem_2_0[0 + 642],mem_2_0[0 + 643],mem_2_0[0 + 644],mem_2_0[0 + 645],mem_2_0[0 + 646],mem_2_0[0 + 647],mem_2_0[0 + 648],mem_2_0[0 + 649],mem_2_0[0 + 650],mem_2_0[0 + 651],mem_2_0[0 + 652],mem_2_0[0 + 653],mem_2_0[0 + 654],mem_2_0[0 + 655],mem_2_0[0 + 656],mem_2_0[0 + 657],mem_2_0[0 + 658],mem_2_0[0 + 659],mem_2_0[0 + 660],mem_2_0[0 + 661],mem_2_0[0 + 662],mem_2_0[0 + 663],mem_2_0[0 + 664],mem_2_0[0 + 665],mem_2_0[0 + 666],mem_2_0[0 + 667],mem_2_0[0 + 668],mem_2_0[0 + 669],mem_2_0[0 + 670],mem_2_0[0 + 671],mem_2_0[0 + 672],mem_2_0[0 + 673],mem_2_0[0 + 674],mem_2_0[0 + 675],mem_2_0[0 + 676],mem_2_0[0 + 677],mem_2_0[0 + 678],mem_2_0[0 + 679],mem_2_0[0 + 680],mem_2_0[0 + 681],mem_2_0[0 + 682],mem_2_0[0 + 683],mem_2_0[0 + 684],mem_2_0[0 + 685],mem_2_0[0 + 686],mem_2_0[0 + 687],mem_2_0[0 + 688],mem_2_0[0 + 689],mem_2_0[0 + 690],mem_2_0[0 + 691],mem_2_0[0 + 692],mem_2_0[0 + 693],mem_2_0[0 + 694],mem_2_0[0 + 695],mem_2_0[0 + 696],mem_2_0[0 + 697],mem_2_0[0 + 698],mem_2_0[0 + 699],mem_2_0[0 + 700],mem_2_0[0 + 701],mem_2_0[0 + 702],mem_2_0[0 + 703],mem_2_0[0 + 704],mem_2_0[0 + 705],mem_2_0[0 + 706],mem_2_0[0 + 707],mem_2_0[0 + 708],mem_2_0[0 + 709],mem_2_0[0 + 710],mem_2_0[0 + 711],mem_2_0[0 + 712],mem_2_0[0 + 713],mem_2_0[0 + 714],mem_2_0[0 + 715],mem_2_0[0 + 716],mem_2_0[0 + 717],mem_2_0[0 + 718],mem_2_0[0 + 719],mem_2_0[0 + 720],mem_2_0[0 + 721],mem_2_0[0 + 722],mem_2_0[0 + 723],mem_2_0[0 + 724],mem_2_0[0 + 725],mem_2_0[0 + 726],mem_2_0[0 + 727],mem_2_0[0 + 728],mem_2_0[0 + 729],mem_2_0[0 + 730],mem_2_0[0 + 731],mem_2_0[0 + 732],mem_2_0[0 + 733],mem_2_0[0 + 734],mem_2_0[0 + 735],mem_2_0[0 + 736],mem_2_0[0 + 737],mem_2_0[0 + 738],mem_2_0[0 + 739],mem_2_0[0 + 740],mem_2_0[0 + 741],mem_2_0[0 + 742],mem_2_0[0 + 743],mem_2_0[0 + 744],mem_2_0[0 + 745],mem_2_0[0 + 746],mem_2_0[0 + 747],mem_2_0[0 + 748],mem_2_0[0 + 749],mem_2_0[0 + 750],mem_2_0[0 + 751],mem_2_0[0 + 752],mem_2_0[0 + 753],mem_2_0[0 + 754],mem_2_0[0 + 755],mem_2_0[0 + 756],mem_2_0[0 + 757],mem_2_0[0 + 758],mem_2_0[0 + 759],mem_2_0[0 + 760],mem_2_0[0 + 761],mem_2_0[0 + 762],mem_2_0[0 + 763],mem_2_0[0 + 764],mem_2_0[0 + 765],mem_2_0[0 + 766],mem_2_0[0 + 767],mem_2_0[0 + 768],mem_2_0[0 + 769],mem_2_0[0 + 770],mem_2_0[0 + 771],mem_2_0[0 + 772],mem_2_0[0 + 773],mem_2_0[0 + 774],mem_2_0[0 + 775],mem_2_0[0 + 776],mem_2_0[0 + 777],mem_2_0[0 + 778],mem_2_0[0 + 779],mem_2_0[0 + 780],mem_2_0[0 + 781],mem_2_0[0 + 782],mem_2_0[0 + 783],mem_2_0[0 + 784],mem_2_0[0 + 785],mem_2_0[0 + 786],mem_2_0[0 + 787],mem_2_0[0 + 788],mem_2_0[0 + 789],mem_2_0[0 + 790],mem_2_0[0 + 791],mem_2_0[0 + 792],mem_2_0[0 + 793],mem_2_0[0 + 794],mem_2_0[0 + 795],mem_2_0[0 + 796],mem_2_0[0 + 797],mem_2_0[0 + 798],mem_2_0[0 + 799],mem_2_0[0 + 800],mem_2_0[0 + 801],mem_2_0[0 + 802],mem_2_0[0 + 803],mem_2_0[0 + 804],mem_2_0[0 + 805],mem_2_0[0 + 806],mem_2_0[0 + 807],mem_2_0[0 + 808],mem_2_0[0 + 809],mem_2_0[0 + 810],mem_2_0[0 + 811],mem_2_0[0 + 812],mem_2_0[0 + 813],mem_2_0[0 + 814],mem_2_0[0 + 815],mem_2_0[0 + 816],mem_2_0[0 + 817],mem_2_0[0 + 818],mem_2_0[0 + 819],mem_2_0[0 + 820],mem_2_0[0 + 821],mem_2_0[0 + 822],mem_2_0[0 + 823],mem_2_0[0 + 824],mem_2_0[0 + 825],mem_2_0[0 + 826],mem_2_0[0 + 827],mem_2_0[0 + 828],mem_2_0[0 + 829],mem_2_0[0 + 830],mem_2_0[0 + 831],mem_2_0[0 + 832],mem_2_0[0 + 833],mem_2_0[0 + 834],mem_2_0[0 + 835],mem_2_0[0 + 836],mem_2_0[0 + 837],mem_2_0[0 + 838],mem_2_0[0 + 839],mem_2_0[0 + 840],mem_2_0[0 + 841],mem_2_0[0 + 842],mem_2_0[0 + 843],mem_2_0[0 + 844],mem_2_0[0 + 845],mem_2_0[0 + 846],mem_2_0[0 + 847],mem_2_0[0 + 848],mem_2_0[0 + 849],mem_2_0[0 + 850],mem_2_0[0 + 851],mem_2_0[0 + 852],mem_2_0[0 + 853],mem_2_0[0 + 854],mem_2_0[0 + 855],mem_2_0[0 + 856],mem_2_0[0 + 857],mem_2_0[0 + 858],mem_2_0[0 + 859],mem_2_0[0 + 860],mem_2_0[0 + 861],mem_2_0[0 + 862],mem_2_0[0 + 863],mem_2_0[0 + 864],mem_2_0[0 + 865],mem_2_0[0 + 866],mem_2_0[0 + 867],mem_2_0[0 + 868],mem_2_0[0 + 869],mem_2_0[0 + 870],mem_2_0[0 + 871],mem_2_0[0 + 872],mem_2_0[0 + 873],mem_2_0[0 + 874],mem_2_0[0 + 875],mem_2_0[0 + 876],mem_2_0[0 + 877],mem_2_0[0 + 878],mem_2_0[0 + 879],mem_2_0[0 + 880],mem_2_0[0 + 881],mem_2_0[0 + 882],mem_2_0[0 + 883],mem_2_0[0 + 884],mem_2_0[0 + 885],mem_2_0[0 + 886],mem_2_0[0 + 887],mem_2_0[0 + 888],mem_2_0[0 + 889],mem_2_0[0 + 890],mem_2_0[0 + 891],mem_2_0[0 + 892],mem_2_0[0 + 893],mem_2_0[0 + 894],mem_2_0[0 + 895],mem_2_0[0 + 896],mem_2_0[0 + 897],mem_2_0[0 + 898],mem_2_0[0 + 899],mem_2_0[0 + 900],mem_2_0[0 + 901],mem_2_0[0 + 902],mem_2_0[0 + 903],mem_2_0[0 + 904],mem_2_0[0 + 905],mem_2_0[0 + 906],mem_2_0[0 + 907],mem_2_0[0 + 908],mem_2_0[0 + 909],mem_2_0[0 + 910],mem_2_0[0 + 911],mem_2_0[0 + 912],mem_2_0[0 + 913],mem_2_0[0 + 914],mem_2_0[0 + 915],mem_2_0[0 + 916],mem_2_0[0 + 917],mem_2_0[0 + 918],mem_2_0[0 + 919],mem_2_0[0 + 920],mem_2_0[0 + 921],mem_2_0[0 + 922],mem_2_0[0 + 923],mem_2_0[0 + 924],mem_2_0[0 + 925],mem_2_0[0 + 926],mem_2_0[0 + 927],mem_2_0[0 + 928],mem_2_0[0 + 929],mem_2_0[0 + 930],mem_2_0[0 + 931],mem_2_0[0 + 932],mem_2_0[0 + 933],mem_2_0[0 + 934],mem_2_0[0 + 935],mem_2_0[0 + 936],mem_2_0[0 + 937],mem_2_0[0 + 938],mem_2_0[0 + 939],mem_2_0[0 + 940],mem_2_0[0 + 941],mem_2_0[0 + 942],mem_2_0[0 + 943],mem_2_0[0 + 944],mem_2_0[0 + 945],mem_2_0[0 + 946],mem_2_0[0 + 947],mem_2_0[0 + 948],mem_2_0[0 + 949],mem_2_0[0 + 950],mem_2_0[0 + 951],mem_2_0[0 + 952],mem_2_0[0 + 953],mem_2_0[0 + 954],mem_2_0[0 + 955],mem_2_0[0 + 956],mem_2_0[0 + 957],mem_2_0[0 + 958],mem_2_0[0 + 959],mem_2_0[0 + 960],mem_2_0[0 + 961],mem_2_0[0 + 962],mem_2_0[0 + 963],mem_2_0[0 + 964],mem_2_0[0 + 965],mem_2_0[0 + 966],mem_2_0[0 + 967],mem_2_0[0 + 968],mem_2_0[0 + 969],mem_2_0[0 + 970],mem_2_0[0 + 971],mem_2_0[0 + 972],mem_2_0[0 + 973],mem_2_0[0 + 974],mem_2_0[0 + 975],mem_2_0[0 + 976],mem_2_0[0 + 977],mem_2_0[0 + 978],mem_2_0[0 + 979],mem_2_0[0 + 980],mem_2_0[0 + 981],mem_2_0[0 + 982],mem_2_0[0 + 983],mem_2_0[0 + 984],mem_2_0[0 + 985],mem_2_0[0 + 986],mem_2_0[0 + 987],mem_2_0[0 + 988],mem_2_0[0 + 989],mem_2_0[0 + 990],mem_2_0[0 + 991],mem_2_0[0 + 992],mem_2_0[0 + 993],mem_2_0[0 + 994],mem_2_0[0 + 995],mem_2_0[0 + 996],mem_2_0[0 + 997],mem_2_0[0 + 998],mem_2_0[0 + 999],mem_2_0[0 + 1000],mem_2_0[0 + 1001],mem_2_0[0 + 1002],mem_2_0[0 + 1003],mem_2_0[0 + 1004],mem_2_0[0 + 1005],mem_2_0[0 + 1006],mem_2_0[0 + 1007],mem_2_0[0 + 1008],mem_2_0[0 + 1009],mem_2_0[0 + 1010],mem_2_0[0 + 1011],mem_2_0[0 + 1012],mem_2_0[0 + 1013],mem_2_0[0 + 1014],mem_2_0[0 + 1015],mem_2_0[0 + 1016],mem_2_0[0 + 1017],mem_2_0[0 + 1018],mem_2_0[0 + 1019],mem_2_0[0 + 1020],mem_2_0[0 + 1021],mem_2_0[0 + 1022],mem_2_0[0 + 1024 - 1] };
wire [8*(1024)-1:0] mem_3_0_flat_src;
assign mem_3_0_flat_src = {mem_3_0[0 + 0],mem_3_0[0 + 1],mem_3_0[0 + 2],mem_3_0[0 + 3],mem_3_0[0 + 4],mem_3_0[0 + 5],mem_3_0[0 + 6],mem_3_0[0 + 7],mem_3_0[0 + 8],mem_3_0[0 + 9],mem_3_0[0 + 10],mem_3_0[0 + 11],mem_3_0[0 + 12],mem_3_0[0 + 13],mem_3_0[0 + 14],mem_3_0[0 + 15],mem_3_0[0 + 16],mem_3_0[0 + 17],mem_3_0[0 + 18],mem_3_0[0 + 19],mem_3_0[0 + 20],mem_3_0[0 + 21],mem_3_0[0 + 22],mem_3_0[0 + 23],mem_3_0[0 + 24],mem_3_0[0 + 25],mem_3_0[0 + 26],mem_3_0[0 + 27],mem_3_0[0 + 28],mem_3_0[0 + 29],mem_3_0[0 + 30],mem_3_0[0 + 31],mem_3_0[0 + 32],mem_3_0[0 + 33],mem_3_0[0 + 34],mem_3_0[0 + 35],mem_3_0[0 + 36],mem_3_0[0 + 37],mem_3_0[0 + 38],mem_3_0[0 + 39],mem_3_0[0 + 40],mem_3_0[0 + 41],mem_3_0[0 + 42],mem_3_0[0 + 43],mem_3_0[0 + 44],mem_3_0[0 + 45],mem_3_0[0 + 46],mem_3_0[0 + 47],mem_3_0[0 + 48],mem_3_0[0 + 49],mem_3_0[0 + 50],mem_3_0[0 + 51],mem_3_0[0 + 52],mem_3_0[0 + 53],mem_3_0[0 + 54],mem_3_0[0 + 55],mem_3_0[0 + 56],mem_3_0[0 + 57],mem_3_0[0 + 58],mem_3_0[0 + 59],mem_3_0[0 + 60],mem_3_0[0 + 61],mem_3_0[0 + 62],mem_3_0[0 + 63],mem_3_0[0 + 64],mem_3_0[0 + 65],mem_3_0[0 + 66],mem_3_0[0 + 67],mem_3_0[0 + 68],mem_3_0[0 + 69],mem_3_0[0 + 70],mem_3_0[0 + 71],mem_3_0[0 + 72],mem_3_0[0 + 73],mem_3_0[0 + 74],mem_3_0[0 + 75],mem_3_0[0 + 76],mem_3_0[0 + 77],mem_3_0[0 + 78],mem_3_0[0 + 79],mem_3_0[0 + 80],mem_3_0[0 + 81],mem_3_0[0 + 82],mem_3_0[0 + 83],mem_3_0[0 + 84],mem_3_0[0 + 85],mem_3_0[0 + 86],mem_3_0[0 + 87],mem_3_0[0 + 88],mem_3_0[0 + 89],mem_3_0[0 + 90],mem_3_0[0 + 91],mem_3_0[0 + 92],mem_3_0[0 + 93],mem_3_0[0 + 94],mem_3_0[0 + 95],mem_3_0[0 + 96],mem_3_0[0 + 97],mem_3_0[0 + 98],mem_3_0[0 + 99],mem_3_0[0 + 100],mem_3_0[0 + 101],mem_3_0[0 + 102],mem_3_0[0 + 103],mem_3_0[0 + 104],mem_3_0[0 + 105],mem_3_0[0 + 106],mem_3_0[0 + 107],mem_3_0[0 + 108],mem_3_0[0 + 109],mem_3_0[0 + 110],mem_3_0[0 + 111],mem_3_0[0 + 112],mem_3_0[0 + 113],mem_3_0[0 + 114],mem_3_0[0 + 115],mem_3_0[0 + 116],mem_3_0[0 + 117],mem_3_0[0 + 118],mem_3_0[0 + 119],mem_3_0[0 + 120],mem_3_0[0 + 121],mem_3_0[0 + 122],mem_3_0[0 + 123],mem_3_0[0 + 124],mem_3_0[0 + 125],mem_3_0[0 + 126],mem_3_0[0 + 127],mem_3_0[0 + 128],mem_3_0[0 + 129],mem_3_0[0 + 130],mem_3_0[0 + 131],mem_3_0[0 + 132],mem_3_0[0 + 133],mem_3_0[0 + 134],mem_3_0[0 + 135],mem_3_0[0 + 136],mem_3_0[0 + 137],mem_3_0[0 + 138],mem_3_0[0 + 139],mem_3_0[0 + 140],mem_3_0[0 + 141],mem_3_0[0 + 142],mem_3_0[0 + 143],mem_3_0[0 + 144],mem_3_0[0 + 145],mem_3_0[0 + 146],mem_3_0[0 + 147],mem_3_0[0 + 148],mem_3_0[0 + 149],mem_3_0[0 + 150],mem_3_0[0 + 151],mem_3_0[0 + 152],mem_3_0[0 + 153],mem_3_0[0 + 154],mem_3_0[0 + 155],mem_3_0[0 + 156],mem_3_0[0 + 157],mem_3_0[0 + 158],mem_3_0[0 + 159],mem_3_0[0 + 160],mem_3_0[0 + 161],mem_3_0[0 + 162],mem_3_0[0 + 163],mem_3_0[0 + 164],mem_3_0[0 + 165],mem_3_0[0 + 166],mem_3_0[0 + 167],mem_3_0[0 + 168],mem_3_0[0 + 169],mem_3_0[0 + 170],mem_3_0[0 + 171],mem_3_0[0 + 172],mem_3_0[0 + 173],mem_3_0[0 + 174],mem_3_0[0 + 175],mem_3_0[0 + 176],mem_3_0[0 + 177],mem_3_0[0 + 178],mem_3_0[0 + 179],mem_3_0[0 + 180],mem_3_0[0 + 181],mem_3_0[0 + 182],mem_3_0[0 + 183],mem_3_0[0 + 184],mem_3_0[0 + 185],mem_3_0[0 + 186],mem_3_0[0 + 187],mem_3_0[0 + 188],mem_3_0[0 + 189],mem_3_0[0 + 190],mem_3_0[0 + 191],mem_3_0[0 + 192],mem_3_0[0 + 193],mem_3_0[0 + 194],mem_3_0[0 + 195],mem_3_0[0 + 196],mem_3_0[0 + 197],mem_3_0[0 + 198],mem_3_0[0 + 199],mem_3_0[0 + 200],mem_3_0[0 + 201],mem_3_0[0 + 202],mem_3_0[0 + 203],mem_3_0[0 + 204],mem_3_0[0 + 205],mem_3_0[0 + 206],mem_3_0[0 + 207],mem_3_0[0 + 208],mem_3_0[0 + 209],mem_3_0[0 + 210],mem_3_0[0 + 211],mem_3_0[0 + 212],mem_3_0[0 + 213],mem_3_0[0 + 214],mem_3_0[0 + 215],mem_3_0[0 + 216],mem_3_0[0 + 217],mem_3_0[0 + 218],mem_3_0[0 + 219],mem_3_0[0 + 220],mem_3_0[0 + 221],mem_3_0[0 + 222],mem_3_0[0 + 223],mem_3_0[0 + 224],mem_3_0[0 + 225],mem_3_0[0 + 226],mem_3_0[0 + 227],mem_3_0[0 + 228],mem_3_0[0 + 229],mem_3_0[0 + 230],mem_3_0[0 + 231],mem_3_0[0 + 232],mem_3_0[0 + 233],mem_3_0[0 + 234],mem_3_0[0 + 235],mem_3_0[0 + 236],mem_3_0[0 + 237],mem_3_0[0 + 238],mem_3_0[0 + 239],mem_3_0[0 + 240],mem_3_0[0 + 241],mem_3_0[0 + 242],mem_3_0[0 + 243],mem_3_0[0 + 244],mem_3_0[0 + 245],mem_3_0[0 + 246],mem_3_0[0 + 247],mem_3_0[0 + 248],mem_3_0[0 + 249],mem_3_0[0 + 250],mem_3_0[0 + 251],mem_3_0[0 + 252],mem_3_0[0 + 253],mem_3_0[0 + 254],mem_3_0[0 + 255],mem_3_0[0 + 256],mem_3_0[0 + 257],mem_3_0[0 + 258],mem_3_0[0 + 259],mem_3_0[0 + 260],mem_3_0[0 + 261],mem_3_0[0 + 262],mem_3_0[0 + 263],mem_3_0[0 + 264],mem_3_0[0 + 265],mem_3_0[0 + 266],mem_3_0[0 + 267],mem_3_0[0 + 268],mem_3_0[0 + 269],mem_3_0[0 + 270],mem_3_0[0 + 271],mem_3_0[0 + 272],mem_3_0[0 + 273],mem_3_0[0 + 274],mem_3_0[0 + 275],mem_3_0[0 + 276],mem_3_0[0 + 277],mem_3_0[0 + 278],mem_3_0[0 + 279],mem_3_0[0 + 280],mem_3_0[0 + 281],mem_3_0[0 + 282],mem_3_0[0 + 283],mem_3_0[0 + 284],mem_3_0[0 + 285],mem_3_0[0 + 286],mem_3_0[0 + 287],mem_3_0[0 + 288],mem_3_0[0 + 289],mem_3_0[0 + 290],mem_3_0[0 + 291],mem_3_0[0 + 292],mem_3_0[0 + 293],mem_3_0[0 + 294],mem_3_0[0 + 295],mem_3_0[0 + 296],mem_3_0[0 + 297],mem_3_0[0 + 298],mem_3_0[0 + 299],mem_3_0[0 + 300],mem_3_0[0 + 301],mem_3_0[0 + 302],mem_3_0[0 + 303],mem_3_0[0 + 304],mem_3_0[0 + 305],mem_3_0[0 + 306],mem_3_0[0 + 307],mem_3_0[0 + 308],mem_3_0[0 + 309],mem_3_0[0 + 310],mem_3_0[0 + 311],mem_3_0[0 + 312],mem_3_0[0 + 313],mem_3_0[0 + 314],mem_3_0[0 + 315],mem_3_0[0 + 316],mem_3_0[0 + 317],mem_3_0[0 + 318],mem_3_0[0 + 319],mem_3_0[0 + 320],mem_3_0[0 + 321],mem_3_0[0 + 322],mem_3_0[0 + 323],mem_3_0[0 + 324],mem_3_0[0 + 325],mem_3_0[0 + 326],mem_3_0[0 + 327],mem_3_0[0 + 328],mem_3_0[0 + 329],mem_3_0[0 + 330],mem_3_0[0 + 331],mem_3_0[0 + 332],mem_3_0[0 + 333],mem_3_0[0 + 334],mem_3_0[0 + 335],mem_3_0[0 + 336],mem_3_0[0 + 337],mem_3_0[0 + 338],mem_3_0[0 + 339],mem_3_0[0 + 340],mem_3_0[0 + 341],mem_3_0[0 + 342],mem_3_0[0 + 343],mem_3_0[0 + 344],mem_3_0[0 + 345],mem_3_0[0 + 346],mem_3_0[0 + 347],mem_3_0[0 + 348],mem_3_0[0 + 349],mem_3_0[0 + 350],mem_3_0[0 + 351],mem_3_0[0 + 352],mem_3_0[0 + 353],mem_3_0[0 + 354],mem_3_0[0 + 355],mem_3_0[0 + 356],mem_3_0[0 + 357],mem_3_0[0 + 358],mem_3_0[0 + 359],mem_3_0[0 + 360],mem_3_0[0 + 361],mem_3_0[0 + 362],mem_3_0[0 + 363],mem_3_0[0 + 364],mem_3_0[0 + 365],mem_3_0[0 + 366],mem_3_0[0 + 367],mem_3_0[0 + 368],mem_3_0[0 + 369],mem_3_0[0 + 370],mem_3_0[0 + 371],mem_3_0[0 + 372],mem_3_0[0 + 373],mem_3_0[0 + 374],mem_3_0[0 + 375],mem_3_0[0 + 376],mem_3_0[0 + 377],mem_3_0[0 + 378],mem_3_0[0 + 379],mem_3_0[0 + 380],mem_3_0[0 + 381],mem_3_0[0 + 382],mem_3_0[0 + 383],mem_3_0[0 + 384],mem_3_0[0 + 385],mem_3_0[0 + 386],mem_3_0[0 + 387],mem_3_0[0 + 388],mem_3_0[0 + 389],mem_3_0[0 + 390],mem_3_0[0 + 391],mem_3_0[0 + 392],mem_3_0[0 + 393],mem_3_0[0 + 394],mem_3_0[0 + 395],mem_3_0[0 + 396],mem_3_0[0 + 397],mem_3_0[0 + 398],mem_3_0[0 + 399],mem_3_0[0 + 400],mem_3_0[0 + 401],mem_3_0[0 + 402],mem_3_0[0 + 403],mem_3_0[0 + 404],mem_3_0[0 + 405],mem_3_0[0 + 406],mem_3_0[0 + 407],mem_3_0[0 + 408],mem_3_0[0 + 409],mem_3_0[0 + 410],mem_3_0[0 + 411],mem_3_0[0 + 412],mem_3_0[0 + 413],mem_3_0[0 + 414],mem_3_0[0 + 415],mem_3_0[0 + 416],mem_3_0[0 + 417],mem_3_0[0 + 418],mem_3_0[0 + 419],mem_3_0[0 + 420],mem_3_0[0 + 421],mem_3_0[0 + 422],mem_3_0[0 + 423],mem_3_0[0 + 424],mem_3_0[0 + 425],mem_3_0[0 + 426],mem_3_0[0 + 427],mem_3_0[0 + 428],mem_3_0[0 + 429],mem_3_0[0 + 430],mem_3_0[0 + 431],mem_3_0[0 + 432],mem_3_0[0 + 433],mem_3_0[0 + 434],mem_3_0[0 + 435],mem_3_0[0 + 436],mem_3_0[0 + 437],mem_3_0[0 + 438],mem_3_0[0 + 439],mem_3_0[0 + 440],mem_3_0[0 + 441],mem_3_0[0 + 442],mem_3_0[0 + 443],mem_3_0[0 + 444],mem_3_0[0 + 445],mem_3_0[0 + 446],mem_3_0[0 + 447],mem_3_0[0 + 448],mem_3_0[0 + 449],mem_3_0[0 + 450],mem_3_0[0 + 451],mem_3_0[0 + 452],mem_3_0[0 + 453],mem_3_0[0 + 454],mem_3_0[0 + 455],mem_3_0[0 + 456],mem_3_0[0 + 457],mem_3_0[0 + 458],mem_3_0[0 + 459],mem_3_0[0 + 460],mem_3_0[0 + 461],mem_3_0[0 + 462],mem_3_0[0 + 463],mem_3_0[0 + 464],mem_3_0[0 + 465],mem_3_0[0 + 466],mem_3_0[0 + 467],mem_3_0[0 + 468],mem_3_0[0 + 469],mem_3_0[0 + 470],mem_3_0[0 + 471],mem_3_0[0 + 472],mem_3_0[0 + 473],mem_3_0[0 + 474],mem_3_0[0 + 475],mem_3_0[0 + 476],mem_3_0[0 + 477],mem_3_0[0 + 478],mem_3_0[0 + 479],mem_3_0[0 + 480],mem_3_0[0 + 481],mem_3_0[0 + 482],mem_3_0[0 + 483],mem_3_0[0 + 484],mem_3_0[0 + 485],mem_3_0[0 + 486],mem_3_0[0 + 487],mem_3_0[0 + 488],mem_3_0[0 + 489],mem_3_0[0 + 490],mem_3_0[0 + 491],mem_3_0[0 + 492],mem_3_0[0 + 493],mem_3_0[0 + 494],mem_3_0[0 + 495],mem_3_0[0 + 496],mem_3_0[0 + 497],mem_3_0[0 + 498],mem_3_0[0 + 499],mem_3_0[0 + 500],mem_3_0[0 + 501],mem_3_0[0 + 502],mem_3_0[0 + 503],mem_3_0[0 + 504],mem_3_0[0 + 505],mem_3_0[0 + 506],mem_3_0[0 + 507],mem_3_0[0 + 508],mem_3_0[0 + 509],mem_3_0[0 + 510],mem_3_0[0 + 511],mem_3_0[0 + 512],mem_3_0[0 + 513],mem_3_0[0 + 514],mem_3_0[0 + 515],mem_3_0[0 + 516],mem_3_0[0 + 517],mem_3_0[0 + 518],mem_3_0[0 + 519],mem_3_0[0 + 520],mem_3_0[0 + 521],mem_3_0[0 + 522],mem_3_0[0 + 523],mem_3_0[0 + 524],mem_3_0[0 + 525],mem_3_0[0 + 526],mem_3_0[0 + 527],mem_3_0[0 + 528],mem_3_0[0 + 529],mem_3_0[0 + 530],mem_3_0[0 + 531],mem_3_0[0 + 532],mem_3_0[0 + 533],mem_3_0[0 + 534],mem_3_0[0 + 535],mem_3_0[0 + 536],mem_3_0[0 + 537],mem_3_0[0 + 538],mem_3_0[0 + 539],mem_3_0[0 + 540],mem_3_0[0 + 541],mem_3_0[0 + 542],mem_3_0[0 + 543],mem_3_0[0 + 544],mem_3_0[0 + 545],mem_3_0[0 + 546],mem_3_0[0 + 547],mem_3_0[0 + 548],mem_3_0[0 + 549],mem_3_0[0 + 550],mem_3_0[0 + 551],mem_3_0[0 + 552],mem_3_0[0 + 553],mem_3_0[0 + 554],mem_3_0[0 + 555],mem_3_0[0 + 556],mem_3_0[0 + 557],mem_3_0[0 + 558],mem_3_0[0 + 559],mem_3_0[0 + 560],mem_3_0[0 + 561],mem_3_0[0 + 562],mem_3_0[0 + 563],mem_3_0[0 + 564],mem_3_0[0 + 565],mem_3_0[0 + 566],mem_3_0[0 + 567],mem_3_0[0 + 568],mem_3_0[0 + 569],mem_3_0[0 + 570],mem_3_0[0 + 571],mem_3_0[0 + 572],mem_3_0[0 + 573],mem_3_0[0 + 574],mem_3_0[0 + 575],mem_3_0[0 + 576],mem_3_0[0 + 577],mem_3_0[0 + 578],mem_3_0[0 + 579],mem_3_0[0 + 580],mem_3_0[0 + 581],mem_3_0[0 + 582],mem_3_0[0 + 583],mem_3_0[0 + 584],mem_3_0[0 + 585],mem_3_0[0 + 586],mem_3_0[0 + 587],mem_3_0[0 + 588],mem_3_0[0 + 589],mem_3_0[0 + 590],mem_3_0[0 + 591],mem_3_0[0 + 592],mem_3_0[0 + 593],mem_3_0[0 + 594],mem_3_0[0 + 595],mem_3_0[0 + 596],mem_3_0[0 + 597],mem_3_0[0 + 598],mem_3_0[0 + 599],mem_3_0[0 + 600],mem_3_0[0 + 601],mem_3_0[0 + 602],mem_3_0[0 + 603],mem_3_0[0 + 604],mem_3_0[0 + 605],mem_3_0[0 + 606],mem_3_0[0 + 607],mem_3_0[0 + 608],mem_3_0[0 + 609],mem_3_0[0 + 610],mem_3_0[0 + 611],mem_3_0[0 + 612],mem_3_0[0 + 613],mem_3_0[0 + 614],mem_3_0[0 + 615],mem_3_0[0 + 616],mem_3_0[0 + 617],mem_3_0[0 + 618],mem_3_0[0 + 619],mem_3_0[0 + 620],mem_3_0[0 + 621],mem_3_0[0 + 622],mem_3_0[0 + 623],mem_3_0[0 + 624],mem_3_0[0 + 625],mem_3_0[0 + 626],mem_3_0[0 + 627],mem_3_0[0 + 628],mem_3_0[0 + 629],mem_3_0[0 + 630],mem_3_0[0 + 631],mem_3_0[0 + 632],mem_3_0[0 + 633],mem_3_0[0 + 634],mem_3_0[0 + 635],mem_3_0[0 + 636],mem_3_0[0 + 637],mem_3_0[0 + 638],mem_3_0[0 + 639],mem_3_0[0 + 640],mem_3_0[0 + 641],mem_3_0[0 + 642],mem_3_0[0 + 643],mem_3_0[0 + 644],mem_3_0[0 + 645],mem_3_0[0 + 646],mem_3_0[0 + 647],mem_3_0[0 + 648],mem_3_0[0 + 649],mem_3_0[0 + 650],mem_3_0[0 + 651],mem_3_0[0 + 652],mem_3_0[0 + 653],mem_3_0[0 + 654],mem_3_0[0 + 655],mem_3_0[0 + 656],mem_3_0[0 + 657],mem_3_0[0 + 658],mem_3_0[0 + 659],mem_3_0[0 + 660],mem_3_0[0 + 661],mem_3_0[0 + 662],mem_3_0[0 + 663],mem_3_0[0 + 664],mem_3_0[0 + 665],mem_3_0[0 + 666],mem_3_0[0 + 667],mem_3_0[0 + 668],mem_3_0[0 + 669],mem_3_0[0 + 670],mem_3_0[0 + 671],mem_3_0[0 + 672],mem_3_0[0 + 673],mem_3_0[0 + 674],mem_3_0[0 + 675],mem_3_0[0 + 676],mem_3_0[0 + 677],mem_3_0[0 + 678],mem_3_0[0 + 679],mem_3_0[0 + 680],mem_3_0[0 + 681],mem_3_0[0 + 682],mem_3_0[0 + 683],mem_3_0[0 + 684],mem_3_0[0 + 685],mem_3_0[0 + 686],mem_3_0[0 + 687],mem_3_0[0 + 688],mem_3_0[0 + 689],mem_3_0[0 + 690],mem_3_0[0 + 691],mem_3_0[0 + 692],mem_3_0[0 + 693],mem_3_0[0 + 694],mem_3_0[0 + 695],mem_3_0[0 + 696],mem_3_0[0 + 697],mem_3_0[0 + 698],mem_3_0[0 + 699],mem_3_0[0 + 700],mem_3_0[0 + 701],mem_3_0[0 + 702],mem_3_0[0 + 703],mem_3_0[0 + 704],mem_3_0[0 + 705],mem_3_0[0 + 706],mem_3_0[0 + 707],mem_3_0[0 + 708],mem_3_0[0 + 709],mem_3_0[0 + 710],mem_3_0[0 + 711],mem_3_0[0 + 712],mem_3_0[0 + 713],mem_3_0[0 + 714],mem_3_0[0 + 715],mem_3_0[0 + 716],mem_3_0[0 + 717],mem_3_0[0 + 718],mem_3_0[0 + 719],mem_3_0[0 + 720],mem_3_0[0 + 721],mem_3_0[0 + 722],mem_3_0[0 + 723],mem_3_0[0 + 724],mem_3_0[0 + 725],mem_3_0[0 + 726],mem_3_0[0 + 727],mem_3_0[0 + 728],mem_3_0[0 + 729],mem_3_0[0 + 730],mem_3_0[0 + 731],mem_3_0[0 + 732],mem_3_0[0 + 733],mem_3_0[0 + 734],mem_3_0[0 + 735],mem_3_0[0 + 736],mem_3_0[0 + 737],mem_3_0[0 + 738],mem_3_0[0 + 739],mem_3_0[0 + 740],mem_3_0[0 + 741],mem_3_0[0 + 742],mem_3_0[0 + 743],mem_3_0[0 + 744],mem_3_0[0 + 745],mem_3_0[0 + 746],mem_3_0[0 + 747],mem_3_0[0 + 748],mem_3_0[0 + 749],mem_3_0[0 + 750],mem_3_0[0 + 751],mem_3_0[0 + 752],mem_3_0[0 + 753],mem_3_0[0 + 754],mem_3_0[0 + 755],mem_3_0[0 + 756],mem_3_0[0 + 757],mem_3_0[0 + 758],mem_3_0[0 + 759],mem_3_0[0 + 760],mem_3_0[0 + 761],mem_3_0[0 + 762],mem_3_0[0 + 763],mem_3_0[0 + 764],mem_3_0[0 + 765],mem_3_0[0 + 766],mem_3_0[0 + 767],mem_3_0[0 + 768],mem_3_0[0 + 769],mem_3_0[0 + 770],mem_3_0[0 + 771],mem_3_0[0 + 772],mem_3_0[0 + 773],mem_3_0[0 + 774],mem_3_0[0 + 775],mem_3_0[0 + 776],mem_3_0[0 + 777],mem_3_0[0 + 778],mem_3_0[0 + 779],mem_3_0[0 + 780],mem_3_0[0 + 781],mem_3_0[0 + 782],mem_3_0[0 + 783],mem_3_0[0 + 784],mem_3_0[0 + 785],mem_3_0[0 + 786],mem_3_0[0 + 787],mem_3_0[0 + 788],mem_3_0[0 + 789],mem_3_0[0 + 790],mem_3_0[0 + 791],mem_3_0[0 + 792],mem_3_0[0 + 793],mem_3_0[0 + 794],mem_3_0[0 + 795],mem_3_0[0 + 796],mem_3_0[0 + 797],mem_3_0[0 + 798],mem_3_0[0 + 799],mem_3_0[0 + 800],mem_3_0[0 + 801],mem_3_0[0 + 802],mem_3_0[0 + 803],mem_3_0[0 + 804],mem_3_0[0 + 805],mem_3_0[0 + 806],mem_3_0[0 + 807],mem_3_0[0 + 808],mem_3_0[0 + 809],mem_3_0[0 + 810],mem_3_0[0 + 811],mem_3_0[0 + 812],mem_3_0[0 + 813],mem_3_0[0 + 814],mem_3_0[0 + 815],mem_3_0[0 + 816],mem_3_0[0 + 817],mem_3_0[0 + 818],mem_3_0[0 + 819],mem_3_0[0 + 820],mem_3_0[0 + 821],mem_3_0[0 + 822],mem_3_0[0 + 823],mem_3_0[0 + 824],mem_3_0[0 + 825],mem_3_0[0 + 826],mem_3_0[0 + 827],mem_3_0[0 + 828],mem_3_0[0 + 829],mem_3_0[0 + 830],mem_3_0[0 + 831],mem_3_0[0 + 832],mem_3_0[0 + 833],mem_3_0[0 + 834],mem_3_0[0 + 835],mem_3_0[0 + 836],mem_3_0[0 + 837],mem_3_0[0 + 838],mem_3_0[0 + 839],mem_3_0[0 + 840],mem_3_0[0 + 841],mem_3_0[0 + 842],mem_3_0[0 + 843],mem_3_0[0 + 844],mem_3_0[0 + 845],mem_3_0[0 + 846],mem_3_0[0 + 847],mem_3_0[0 + 848],mem_3_0[0 + 849],mem_3_0[0 + 850],mem_3_0[0 + 851],mem_3_0[0 + 852],mem_3_0[0 + 853],mem_3_0[0 + 854],mem_3_0[0 + 855],mem_3_0[0 + 856],mem_3_0[0 + 857],mem_3_0[0 + 858],mem_3_0[0 + 859],mem_3_0[0 + 860],mem_3_0[0 + 861],mem_3_0[0 + 862],mem_3_0[0 + 863],mem_3_0[0 + 864],mem_3_0[0 + 865],mem_3_0[0 + 866],mem_3_0[0 + 867],mem_3_0[0 + 868],mem_3_0[0 + 869],mem_3_0[0 + 870],mem_3_0[0 + 871],mem_3_0[0 + 872],mem_3_0[0 + 873],mem_3_0[0 + 874],mem_3_0[0 + 875],mem_3_0[0 + 876],mem_3_0[0 + 877],mem_3_0[0 + 878],mem_3_0[0 + 879],mem_3_0[0 + 880],mem_3_0[0 + 881],mem_3_0[0 + 882],mem_3_0[0 + 883],mem_3_0[0 + 884],mem_3_0[0 + 885],mem_3_0[0 + 886],mem_3_0[0 + 887],mem_3_0[0 + 888],mem_3_0[0 + 889],mem_3_0[0 + 890],mem_3_0[0 + 891],mem_3_0[0 + 892],mem_3_0[0 + 893],mem_3_0[0 + 894],mem_3_0[0 + 895],mem_3_0[0 + 896],mem_3_0[0 + 897],mem_3_0[0 + 898],mem_3_0[0 + 899],mem_3_0[0 + 900],mem_3_0[0 + 901],mem_3_0[0 + 902],mem_3_0[0 + 903],mem_3_0[0 + 904],mem_3_0[0 + 905],mem_3_0[0 + 906],mem_3_0[0 + 907],mem_3_0[0 + 908],mem_3_0[0 + 909],mem_3_0[0 + 910],mem_3_0[0 + 911],mem_3_0[0 + 912],mem_3_0[0 + 913],mem_3_0[0 + 914],mem_3_0[0 + 915],mem_3_0[0 + 916],mem_3_0[0 + 917],mem_3_0[0 + 918],mem_3_0[0 + 919],mem_3_0[0 + 920],mem_3_0[0 + 921],mem_3_0[0 + 922],mem_3_0[0 + 923],mem_3_0[0 + 924],mem_3_0[0 + 925],mem_3_0[0 + 926],mem_3_0[0 + 927],mem_3_0[0 + 928],mem_3_0[0 + 929],mem_3_0[0 + 930],mem_3_0[0 + 931],mem_3_0[0 + 932],mem_3_0[0 + 933],mem_3_0[0 + 934],mem_3_0[0 + 935],mem_3_0[0 + 936],mem_3_0[0 + 937],mem_3_0[0 + 938],mem_3_0[0 + 939],mem_3_0[0 + 940],mem_3_0[0 + 941],mem_3_0[0 + 942],mem_3_0[0 + 943],mem_3_0[0 + 944],mem_3_0[0 + 945],mem_3_0[0 + 946],mem_3_0[0 + 947],mem_3_0[0 + 948],mem_3_0[0 + 949],mem_3_0[0 + 950],mem_3_0[0 + 951],mem_3_0[0 + 952],mem_3_0[0 + 953],mem_3_0[0 + 954],mem_3_0[0 + 955],mem_3_0[0 + 956],mem_3_0[0 + 957],mem_3_0[0 + 958],mem_3_0[0 + 959],mem_3_0[0 + 960],mem_3_0[0 + 961],mem_3_0[0 + 962],mem_3_0[0 + 963],mem_3_0[0 + 964],mem_3_0[0 + 965],mem_3_0[0 + 966],mem_3_0[0 + 967],mem_3_0[0 + 968],mem_3_0[0 + 969],mem_3_0[0 + 970],mem_3_0[0 + 971],mem_3_0[0 + 972],mem_3_0[0 + 973],mem_3_0[0 + 974],mem_3_0[0 + 975],mem_3_0[0 + 976],mem_3_0[0 + 977],mem_3_0[0 + 978],mem_3_0[0 + 979],mem_3_0[0 + 980],mem_3_0[0 + 981],mem_3_0[0 + 982],mem_3_0[0 + 983],mem_3_0[0 + 984],mem_3_0[0 + 985],mem_3_0[0 + 986],mem_3_0[0 + 987],mem_3_0[0 + 988],mem_3_0[0 + 989],mem_3_0[0 + 990],mem_3_0[0 + 991],mem_3_0[0 + 992],mem_3_0[0 + 993],mem_3_0[0 + 994],mem_3_0[0 + 995],mem_3_0[0 + 996],mem_3_0[0 + 997],mem_3_0[0 + 998],mem_3_0[0 + 999],mem_3_0[0 + 1000],mem_3_0[0 + 1001],mem_3_0[0 + 1002],mem_3_0[0 + 1003],mem_3_0[0 + 1004],mem_3_0[0 + 1005],mem_3_0[0 + 1006],mem_3_0[0 + 1007],mem_3_0[0 + 1008],mem_3_0[0 + 1009],mem_3_0[0 + 1010],mem_3_0[0 + 1011],mem_3_0[0 + 1012],mem_3_0[0 + 1013],mem_3_0[0 + 1014],mem_3_0[0 + 1015],mem_3_0[0 + 1016],mem_3_0[0 + 1017],mem_3_0[0 + 1018],mem_3_0[0 + 1019],mem_3_0[0 + 1020],mem_3_0[0 + 1021],mem_3_0[0 + 1022],mem_3_0[0 + 1024 - 1] };
endmodule







