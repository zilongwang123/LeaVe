module SodorInternalTile_2stage_invariant ( input [31:0] \Core_2stage.DatPath_2stage.io_imem_resp_bits_data_state_invariant , input [31:0] \Core_2stage.DatPath_2stage.exe_reg_pc , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_eret , input [31:0] \Core_2stage.DatPath_2stage.if_reg_pc , input \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupt , input [31:0] \Core_2stage.DatPath_2stage.io_imem_resp_bits_data , input \Core_2stage.CtlPath_2stage.io_ctl_exception , input \Core_2stage.DatPath_2stage.if_inst_buffer_valid , input \Core_2stage.DatPath_2stage.io_ctl_if_kill_r , input [31:0] \Core_2stage.DatPath_2stage.exe_reg_inst , output io_ctl_exception_invariant_arg0 , output RV32I_invariant_arg0 , output io_eret_invariant_cond , output IF_REG_PC2_invariant_arg0 , output NO_DEFAULT_INST_invariant_arg0 , output NO_DEFAULT_INST_invariant_cond , output IF_INST_BUFFER_VALID_invariant_arg0 , output IF_REG_PC1_invariant_cond , output IF_REG_PC2_invariant_cond , output IF_INST_BUFFER_VALID_invariant_cond , output io_eret_invariant_arg0 , output EXE_REG_PC1_invariant_cond , output io_interrupt_invariant_arg0 , output EXE_REG_PC2_invariant_cond , output io_ctl_exception_invariant_cond , output EXE_REG_INST_invariant_arg0 , output EXE_REG_PC2_invariant_arg0 , output IF_REG_PC1_invariant_arg0 , output io_interrupt_invariant_cond , output RV32I_invariant_cond , output EXE_REG_PC1_invariant_arg0 , output EXE_REG_INST_invariant_cond );
	assign NO_DEFAULT_INST_invariant_cond = 1 ;
	assign NO_DEFAULT_INST_invariant_arg0 = ( ( \Core_2stage.DatPath_2stage.io_imem_resp_bits_data == 32'h4033 ) == 0 ) ;
	assign EXE_REG_INST_invariant_cond = 1 ;
	assign EXE_REG_INST_invariant_arg0 = ( ( \Core_2stage.DatPath_2stage.io_ctl_if_kill_r ) || ( \Core_2stage.DatPath_2stage.exe_reg_inst == \Core_2stage.DatPath_2stage.io_imem_resp_bits_data_state_invariant ) ) ;
	assign EXE_REG_PC1_invariant_cond = 1 ;
	assign EXE_REG_PC1_invariant_arg0 = ( \Core_2stage.DatPath_2stage.exe_reg_pc [1:0] == 0 ) ;
	assign EXE_REG_PC2_invariant_cond = 1 ;
	assign EXE_REG_PC2_invariant_arg0 = ( ( ! \Core_2stage.DatPath_2stage.io_ctl_if_kill_r ) || ( \Core_2stage.DatPath_2stage.exe_reg_pc == 32'h0 ) ) ;
	assign IF_REG_PC1_invariant_cond = 1 ;
	assign IF_REG_PC1_invariant_arg0 =  ( \Core_2stage.DatPath_2stage.if_reg_pc [1:0] == 0 ) ;
	assign IF_REG_PC2_invariant_cond = 1 ;
	assign IF_REG_PC2_invariant_arg0 =  ( ( \Core_2stage.DatPath_2stage.io_ctl_if_kill_r ) || ( \Core_2stage.DatPath_2stage.if_reg_pc == \Core_2stage.DatPath_2stage.exe_reg_pc + 32'h4 ) ) ;
	assign IF_INST_BUFFER_VALID_invariant_cond = 1 ;
	assign IF_INST_BUFFER_VALID_invariant_arg0 =  ( \Core_2stage.DatPath_2stage.if_inst_buffer_valid == 0 ) ;
	assign RV32I_invariant_cond = 1 ;
	assign RV32I_invariant_arg0 =  ( (\Core_2stage.DatPath_2stage.exe_reg_inst [6:0] == 7'h37 ) || (\Core_2stage.DatPath_2stage.exe_reg_inst [6:0] == 7'h17 ) || (\Core_2stage.DatPath_2stage.exe_reg_inst [6:0] == 7'h6f ) || (\Core_2stage.DatPath_2stage.exe_reg_inst [6:0] == 7'h67 ) ||(\Core_2stage.DatPath_2stage.exe_reg_inst [6:0] == 7'h63 ) || (\Core_2stage.DatPath_2stage.exe_reg_inst [6:0] == 7'h3 ) || (\Core_2stage.DatPath_2stage.exe_reg_inst [6:0] == 7'h23 ) || (\Core_2stage.DatPath_2stage.exe_reg_inst [6:0] == 7'h13 ) || (\Core_2stage.DatPath_2stage.exe_reg_inst [6:0] == 7'h33 && (\Core_2stage.DatPath_2stage.exe_reg_inst [31:25] == 7'h0 || \Core_2stage.DatPath_2stage.exe_reg_inst [31:25] == 7'h20 ) ) ) ;
	assign io_ctl_exception_invariant_cond = 1 ;
	assign io_ctl_exception_invariant_arg0 =  ( \Core_2stage.CtlPath_2stage.io_ctl_exception == 0 ) ;
	assign io_eret_invariant_cond = 1 ;
	assign io_eret_invariant_arg0 =  ( \Core_2stage.DatPath_2stage.CSRFile_2stage.io_eret == 0 ) ;
	assign io_interrupt_invariant_cond = 1 ;
	assign io_interrupt_invariant_arg0 =  ( \Core_2stage.DatPath_2stage.CSRFile_2stage.io_interrupt == 0 ) ;
endmodule